PK
     ��/Z.��\n) n)    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_0":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_1":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_2":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_2":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_3":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_4":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_5":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_5":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_6":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_7":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_7":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9":["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_9":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10":["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_10":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_15":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_16":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_17":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_17":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_18":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_18":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_19":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_19":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_20":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_21":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_24":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_24":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_25":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos"],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_29":[],"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_29":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_1_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_1_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_2_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_2_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_2_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_2_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_3_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_3_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_4_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_4_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_5_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_5_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_5_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_5_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_6_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_6_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_6_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_6_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_7_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_7_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_9_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_9_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_10_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_10_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_11_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_11_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_12_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_12_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_12_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_12_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_13_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_13_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos":["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg":["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_16_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_16_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_17_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_17_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_17_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_17_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_18_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_18_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_18_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_18_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_19_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_19_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_19_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_19_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_20_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_20_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_21_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_21_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_22_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_22_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_23_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_23_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_24_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_24_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_24_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_24_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_25_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_25_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_25_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_25_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_26_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_26_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_26_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_26_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_27_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_27_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-neg":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos":["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg":["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4"],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-pos":[],"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg":[],"pin-type-component_150f7ff8-79d3-4bfa-9f54-059e037d3db1_0":[],"pin-type-component_150f7ff8-79d3-4bfa-9f54-059e037d3db1_1":[],"pin-type-component_d1ef43e3-b043-4b2a-bbe7-f2952ece9282_0":[],"pin-type-component_d1ef43e3-b043-4b2a-bbe7-f2952ece9282_1":[],"pin-type-component_39519189-daa3-42d9-a482-f20abb45fb62_0":[],"pin-type-component_39519189-daa3-42d9-a482-f20abb45fb62_1":[],"pin-type-component_81f615f8-ec40-4b71-aed6-27ebc76da0e8_0":[],"pin-type-component_81f615f8-ec40-4b71-aed6-27ebc76da0e8_1":[],"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0"],"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1"],"pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_0":[],"pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_1":[],"pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_2":[],"pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_3":[],"pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_4":[],"pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_5":[],"pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_6":[],"pin-type-component_4d26be02-7540-4873-be49-92b26c548165_0":[],"pin-type-component_4d26be02-7540-4873-be49-92b26c548165_1":[],"pin-type-component_4d26be02-7540-4873-be49-92b26c548165_2":[],"pin-type-component_4d26be02-7540-4873-be49-92b26c548165_3":[],"pin-type-component_4d26be02-7540-4873-be49-92b26c548165_4":[],"pin-type-component_4d26be02-7540-4873-be49-92b26c548165_5":[],"pin-type-component_4d26be02-7540-4873-be49-92b26c548165_6":[],"pin-type-component_4d26be02-7540-4873-be49-92b26c548165_7":[],"pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_0":[],"pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_1":[],"pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_2":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_0":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_1":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_2":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_3":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_4":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_5":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_6":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_7":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_8":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_9":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_10":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_11":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_12":[],"pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_13":[],"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0":["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0"],"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1":["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1"],"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9"],"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos"],"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg"],"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_5":[],"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_6":[],"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_7":[],"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0":["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0"],"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1":["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1"],"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10"],"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos"],"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg"],"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_5":[],"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_6":[],"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_7":[]},"pin_to_color":{"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0":"#189AB4","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_0":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1":"#FF0000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_1":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_2":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_2":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3":"#683D3B","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_3":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4":"#968AE8","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_4":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_5":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_5":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6":"#FF74A3","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_6":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_7":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_7":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8":"#FF0000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8":"#189AB4","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9":"#FFA6FE","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_9":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10":"#774D00","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_10":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11":"#01FFFE","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12":"#968AE8","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12":"#00AE7E","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13":"#FF74A3","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13":"#A75740","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14":"#683D3B","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14":"#98FF52","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_15":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16":"#98FF52","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_16":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_17":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_17":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_18":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_18":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_19":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_19":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20":"#A75740","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_20":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21":"#00AE7E","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_21":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22":"#189AB4","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22":"#01FFFE","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23":"#FF0000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23":"#01FFFE","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_24":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_24":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25":"#FE8900","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_25":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26":"#FE8900","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26":"#FE8900","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27":"#FF0000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28":"#FF0000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_29":"#000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_29":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg":"#189AB4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg":"#189AB4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos":"#FF0000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_1_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_1_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_2_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_2_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_2_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_2_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_3_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_3_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_4_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_4_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_5_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_5_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_5_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_5_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_6_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_6_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_6_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_6_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg":"#189AB4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_7_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_7_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos":"#FF0000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_9_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_9_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_10_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_10_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_11_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_11_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_12_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_12_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_12_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_12_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_13_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_13_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos":"#FF0000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg":"#189AB4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_16_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_16_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_17_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_17_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_17_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_17_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_18_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_18_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_18_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_18_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_19_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_19_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_19_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_19_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_20_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_20_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_21_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_21_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg":"#189AB4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_22_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_22_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos":"#FF0000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_23_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_23_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_24_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_24_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_24_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_24_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_25_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_25_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_25_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_25_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_26_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_26_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_26_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_26_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos":"#FF0000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_27_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_27_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos":"#FF0000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-neg":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos":"#FF0000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg":"#189AB4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-pos":"#000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg":"#000000","pin-type-component_150f7ff8-79d3-4bfa-9f54-059e037d3db1_0":"#000000","pin-type-component_150f7ff8-79d3-4bfa-9f54-059e037d3db1_1":"#000000","pin-type-component_d1ef43e3-b043-4b2a-bbe7-f2952ece9282_0":"#000000","pin-type-component_d1ef43e3-b043-4b2a-bbe7-f2952ece9282_1":"#000000","pin-type-component_39519189-daa3-42d9-a482-f20abb45fb62_0":"#000000","pin-type-component_39519189-daa3-42d9-a482-f20abb45fb62_1":"#000000","pin-type-component_81f615f8-ec40-4b71-aed6-27ebc76da0e8_0":"#000000","pin-type-component_81f615f8-ec40-4b71-aed6-27ebc76da0e8_1":"#000000","pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0":"#FF0000","pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1":"#189AB4","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_0":"#000000","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_1":"#000000","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_2":"#000000","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_3":"#000000","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_4":"#000000","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_5":"#000000","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_6":"#000000","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_0":"#000000","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_1":"#000000","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_2":"#000000","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_3":"#000000","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_4":"#000000","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_5":"#000000","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_6":"#000000","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_7":"#000000","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_0":"#000000","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_1":"#000000","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_2":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_0":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_1":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_2":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_3":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_4":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_5":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_6":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_7":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_8":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_9":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_10":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_11":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_12":"#000000","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_13":"#000000","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0":"#FF0000","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1":"#189AB4","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2":"#FFA6FE","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3":"#FF0000","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4":"#189AB4","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_5":"#000000","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_6":"#000000","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_7":"#000000","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0":"#FF0000","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1":"#189AB4","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2":"#774D00","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3":"#FF0000","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4":"#189AB4","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_5":"#000000","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_6":"#000000","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_7":"#000000"},"pin_to_state":{"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_0":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_1":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_2":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_2":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_3":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_4":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_5":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_5":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_6":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_7":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_7":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_9":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_10":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_15":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_16":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_17":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_17":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_18":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_18":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_19":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_19":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_20":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_21":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_24":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_24":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_25":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_29":"neutral","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_29":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_1_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_1_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_2_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_2_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_2_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_2_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_3_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_3_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_4_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_4_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_5_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_5_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_5_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_5_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_6_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_6_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_6_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_6_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_7_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_7_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_9_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_9_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_10_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_10_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_11_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_11_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_12_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_12_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_12_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_12_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_13_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_13_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_16_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_16_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_17_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_17_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_17_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_17_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_18_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_18_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_18_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_18_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_19_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_19_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_19_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_19_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_20_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_20_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_21_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_21_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_22_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_22_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_23_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_23_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_24_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_24_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_24_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_24_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_25_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_25_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_25_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_25_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_26_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_26_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_26_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_26_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_27_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_27_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-pos":"neutral","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg":"neutral","pin-type-component_150f7ff8-79d3-4bfa-9f54-059e037d3db1_0":"neutral","pin-type-component_150f7ff8-79d3-4bfa-9f54-059e037d3db1_1":"neutral","pin-type-component_d1ef43e3-b043-4b2a-bbe7-f2952ece9282_0":"neutral","pin-type-component_d1ef43e3-b043-4b2a-bbe7-f2952ece9282_1":"neutral","pin-type-component_39519189-daa3-42d9-a482-f20abb45fb62_0":"neutral","pin-type-component_39519189-daa3-42d9-a482-f20abb45fb62_1":"neutral","pin-type-component_81f615f8-ec40-4b71-aed6-27ebc76da0e8_0":"neutral","pin-type-component_81f615f8-ec40-4b71-aed6-27ebc76da0e8_1":"neutral","pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0":"neutral","pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1":"neutral","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_0":"neutral","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_1":"neutral","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_2":"neutral","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_3":"neutral","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_4":"neutral","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_5":"neutral","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_6":"neutral","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_0":"neutral","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_1":"neutral","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_2":"neutral","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_3":"neutral","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_4":"neutral","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_5":"neutral","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_6":"neutral","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_7":"neutral","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_0":"neutral","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_1":"neutral","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_2":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_0":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_1":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_2":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_3":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_4":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_5":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_6":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_7":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_8":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_9":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_10":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_11":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_12":"neutral","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_13":"neutral","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0":"neutral","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1":"neutral","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2":"neutral","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3":"neutral","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4":"neutral","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_5":"neutral","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_6":"neutral","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_7":"neutral","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0":"neutral","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1":"neutral","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2":"neutral","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3":"neutral","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4":"neutral","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_5":"neutral","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_6":"neutral","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_7":"neutral"},"next_color_idx":29,"wires_placed_in_order":[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_0","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-neg"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-pos"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28"],["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-pos"],["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-neg"],["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-neg"],["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-neg"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_16","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-neg","pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_0"],["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-pos"],["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-neg"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-neg","pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9","pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_2"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10","pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_2"],["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_2","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9"],["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_2","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-pos","pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_10"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-neg","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-neg"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos"],["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-neg"],["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11"],["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10"],["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0"],["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3"],["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"],["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1"],["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-pos"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2"],["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_0","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_0","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-neg"]],[]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8"]]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg"]]],[[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg"]],[]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-pos"]]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]],[]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-pos"]]],[[],[["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-neg"]]],[[],[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-neg"]]],[[],[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-pos"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-neg"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-neg"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos"]]],[[["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-pos"]],[]],[[["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-neg"]],[]],[[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-pos"]],[]],[[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-neg"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_16","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_16","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_15","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-neg","pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_0"]]],[[],[["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-pos"]]],[[],[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-neg"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-neg","pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9","pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_2"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10","pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_2"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10","pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_2"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9","pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_2"]],[]],[[],[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_2","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9"]]],[[],[["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_2","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10"]]],[[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-neg"]],[]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-pos","pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_10"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_10","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-neg","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-neg"]]],[[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-neg","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-neg"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26"]]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg"]],[]],[[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-pos"]],[]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg"]]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos"]]],[[],[]],[[],[]],[[["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-neg"]],[]],[[["pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-pos"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10","pin-type-component_cbd318ac-cd25-4f7a-ab31-677022121b06_2"]],[]],[[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-neg"]],[]],[[["pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-pos"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9","pin-type-component_242ef558-8a6d-4765-86dd-ba97e80a9f30_2"]],[]],[[],[["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-neg"]]],[[],[["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11"]]],[[],[["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10"]]],[[["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-neg"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2"]],[]],[[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2"]],[]],[[],[["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0"]]],[[],[["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1"]]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"]]],[[["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"]],[]],[[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"]],[]],[[["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0"]],[]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"]]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3"]]],[[],[["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4"]]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0"]]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0"]]],[[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"]],[]],[[["pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1","pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1"]],[]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1"]]],[[],[["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1"]]],[[],[["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-pos"]]],[[["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-pos"]],[]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2"]]],[[],[["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0":"0000000000000002","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_0":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1":"0000000000000001","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_1":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_2":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_2":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3":"0000000000000011","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_3":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4":"0000000000000010","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_4":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_5":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_5":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6":"0000000000000012","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_6":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_7":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_7":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8":"0000000000000000","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8":"0000000000000003","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9":"0000000000000015","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_9":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10":"0000000000000016","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_10":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_11":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11":"0000000000000023","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12":"0000000000000010","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12":"0000000000000020","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13":"0000000000000012","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13":"0000000000000021","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14":"0000000000000011","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14":"0000000000000019","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_15":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_15":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16":"0000000000000019","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_16":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_17":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_17":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_18":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_18":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_19":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_19":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20":"0000000000000021","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_20":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21":"0000000000000020","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_21":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22":"0000000000000009","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22":"0000000000000023","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23":"0000000000000008","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23":"0000000000000023","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_24":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_24":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25":"0000000000000022","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_25":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26":"0000000000000022","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26":"0000000000000022","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_27":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27":"0000000000000004","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_28":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28":"0000000000000007","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_29":"_","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_29":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg":"0000000000000002","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg":"0000000000000002","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos":"0000000000000001","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_1_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_1_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_2_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_2_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_2_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_2_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_3_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_3_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_3_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_4_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_4_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_4_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_5_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_5_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_5_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_5_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_6_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_6_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_6_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_6_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg":"0000000000000003","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_7_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_7_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos":"0000000000000000","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_8_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_9_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_9_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_9_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_10_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_10_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_10_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_11_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_11_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_11_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_12_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_12_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_12_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_12_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_13_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_13_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_13_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_14_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos":"0000000000000006","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_15_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg":"0000000000000005","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_16_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_16_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_16_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_17_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_17_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_17_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_17_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_18_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_18_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_18_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_18_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_19_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_19_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_19_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_19_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_20_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_20_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_20_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_21_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_21_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_21_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg":"0000000000000009","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_22_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_22_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos":"0000000000000008","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_23_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_23_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_24_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_24_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_24_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_24_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_25_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_25_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_25_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_25_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_26_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_26_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_26_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_26_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos":"0000000000000004","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_27_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_27_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_28_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos":"0000000000000007","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-neg":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos":"0000000000000013","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg":"0000000000000014","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-pos":"_","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_29_polarity-neg":"_","pin-type-component_150f7ff8-79d3-4bfa-9f54-059e037d3db1_0":"_","pin-type-component_150f7ff8-79d3-4bfa-9f54-059e037d3db1_1":"_","pin-type-component_d1ef43e3-b043-4b2a-bbe7-f2952ece9282_0":"_","pin-type-component_d1ef43e3-b043-4b2a-bbe7-f2952ece9282_1":"_","pin-type-component_39519189-daa3-42d9-a482-f20abb45fb62_0":"_","pin-type-component_39519189-daa3-42d9-a482-f20abb45fb62_1":"_","pin-type-component_81f615f8-ec40-4b71-aed6-27ebc76da0e8_0":"_","pin-type-component_81f615f8-ec40-4b71-aed6-27ebc76da0e8_1":"_","pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0":"0000000000000006","pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1":"0000000000000005","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_0":"_","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_1":"_","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_2":"_","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_3":"_","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_4":"_","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_5":"_","pin-type-component_3e0c97b1-8b73-4276-87c5-f4908c2761cb_6":"_","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_0":"_","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_1":"_","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_2":"_","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_3":"_","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_4":"_","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_5":"_","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_6":"_","pin-type-component_4d26be02-7540-4873-be49-92b26c548165_7":"_","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_0":"_","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_1":"_","pin-type-component_143e3a33-8438-4b9b-a254-a1d18f1c065a_2":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_0":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_1":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_2":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_3":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_4":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_5":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_6":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_7":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_8":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_9":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_10":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_11":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_12":"_","pin-type-component_2b1e4dc7-7a05-4105-b1c2-0ed5598fd491_13":"_","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0":"0000000000000006","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1":"0000000000000005","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2":"0000000000000015","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3":"0000000000000013","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4":"0000000000000014","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_5":"_","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_6":"_","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_7":"_","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0":"0000000000000006","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1":"0000000000000005","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2":"0000000000000016","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3":"0000000000000013","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4":"0000000000000014","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_5":"_","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_6":"_","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_7":"_"},"component_id_to_pins":{"150f7ff8-79d3-4bfa-9f54-059e037d3db1":["0","1"],"d1ef43e3-b043-4b2a-bbe7-f2952ece9282":["0","1"],"39519189-daa3-42d9-a482-f20abb45fb62":["0","1"],"81f615f8-ec40-4b71-aed6-27ebc76da0e8":["0","1"],"a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9":["0","1"],"3e0c97b1-8b73-4276-87c5-f4908c2761cb":["0","1","2","3","4","5","6"],"4d26be02-7540-4873-be49-92b26c548165":["0","1","2","3","4","5","6","7"],"143e3a33-8438-4b9b-a254-a1d18f1c065a":["0","1","2"],"2b1e4dc7-7a05-4105-b1c2-0ed5598fd491":["0","1","2","3","4","5","6","7","8","9","10","11","12","13"],"e856bf6f-239f-495d-9f01-2780e496b019":["0","1","2","3","4","5","6","7"],"846761e3-79a5-45ce-9f89-d8258e1f2e70":["0","1","2","3","4","5","6","7"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos"],"0000000000000001":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos"],"0000000000000002":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg"],"0000000000000003":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8"],"0000000000000008":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23"],"0000000000000009":["pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22"],"0000000000000020":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21"],"0000000000000011":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14"],"0000000000000012":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13"],"0000000000000010":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4"],"0000000000000019":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16"],"0000000000000021":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20"],"0000000000000023":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23"],"0000000000000022":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26","pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26"],"0000000000000004":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos"],"0000000000000007":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos"],"0000000000000005":["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1"],"0000000000000006":["pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0"],"0000000000000013":["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3"],"0000000000000014":["pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4","pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4"],"0000000000000015":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9","pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2"],"0000000000000016":["pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10","pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000020":"Net 20","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000010":"Net 10","0000000000000019":"Net 19","0000000000000021":"Net 21","0000000000000023":"Net 23","0000000000000022":"Net 22","0000000000000004":"Net 4","0000000000000007":"Net 7","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16"},"all_breadboard_info_list":["a818362a-9609-419e-afdb-0484a3ad4904_30_2_True_1060_340_up"],"breadboard_info_list":["a818362a-9609-419e-afdb-0484a3ad4904_30_2_True_1060_340_up"],"componentsData":[{"compProperties":{},"position":[1474.4253985,565.882505],"typeId":"2f403b15-90c3-4075-86a3-7ea6b108dda1","componentVersion":1,"instanceId":"a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9","orientation":"left","circleData":[[1367.5,560],[1367.5,575]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"75000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"4","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[1210.0000000000002,695],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"150f7ff8-79d3-4bfa-9f54-059e037d3db1","orientation":"up","circleData":[[1172.5,695],[1247.5000000000005,695]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"100000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"4","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[1203.5721189654346,680],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"39519189-daa3-42d9-a482-f20abb45fb62","orientation":"up","circleData":[[1172.5,680],[1232.5,680]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1181.2503370000004,395.92027400000006],"typeId":"cc6ddea1-99fb-411d-bfec-02f29cfc7b20","componentVersion":3,"instanceId":"3e0c97b1-8b73-4276-87c5-f4908c2761cb","orientation":"up","circleData":[[1067.5,350],[1067.5,365.00000000000006],[1067.5,380.00000000000006],[1067.5,394.99999999999994],[1067.5,410],[1067.5,424.99999999999994],[1067.5,440.00000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[998.9588229999997,642.420944],"typeId":"70f88287-3db7-454f-a714-3fcb737f1bfe","componentVersion":1,"instanceId":"4d26be02-7540-4873-be49-92b26c548165","orientation":"right","circleData":[[1037.5,590],[1037.5,605],[1037.5,620],[1037.5,635],[1037.5,650],[1037.5,665],[1037.5,680],[1037.5,695]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Type":{"version":2,"id":"Type","label":"Type","description":"","units":"","type":"string","value":"LM317","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Type","unit":"","userVisible":true,"required":true}},"position":[1204.2377499999998,754.2469999999998],"typeId":"0a0aa907-9846-42ff-9576-36638174fe13","componentVersion":1,"instanceId":"143e3a33-8438-4b9b-a254-a1d18f1c065a","orientation":"right","circleData":[[1142.5,740],[1142.5,754.997],[1142.5,769.9939999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"330","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"4","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[999.5714745976957,725],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"d1ef43e3-b043-4b2a-bbe7-f2952ece9282","orientation":"up","circleData":[[962.5000000000002,725],[1037.4999999999998,725]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"1000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"4","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[1006.8580173562168,740],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"81f615f8-ec40-4b71-aed6-27ebc76da0e8","orientation":"up","circleData":[[977.5000000000002,740],[1037.5000000000005,740]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1105.0391815,514.649396],"typeId":"7799e1c0-2491-44a2-a64d-b6a1e1bb7939","componentVersion":2,"instanceId":"2b1e4dc7-7a05-4105-b1c2-0ed5598fd491","orientation":"up","circleData":[[1082.5,470],[1082.5,485],[1082.5,500],[1082.5,515],[1082.5,530],[1082.5,545],[1082.5,560],[1127.5,560],[1127.5,545],[1127.5,530],[1127.5,515],[1127.5,500],[1127.5,485],[1127.5,470]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[681.7754605000005,1045.8981650000005],"typeId":"e60aba2b-e9b2-4ddc-8d1b-286ba98ca1ae","componentVersion":1,"instanceId":"846761e3-79a5-45ce-9f89-d8258e1f2e70","orientation":"down","circleData":[[812.5,1009.9999999999998],[813.4210525000003,1073.5526314999997],[845.8690314999998,1049.4629345000003],[833.623099,1042.8358475],[847.951336,1035.1584185000002],[525.717271,1070.3736064999998],[525.717271,1041.9534470000003],[523.9985769999997,1013.5949945]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[681.7754605000002,910.8981650000001],"typeId":"e60aba2b-e9b2-4ddc-8d1b-286ba98ca1ae","componentVersion":1,"instanceId":"e856bf6f-239f-495d-9f01-2780e496b019","orientation":"down","circleData":[[812.5,875],[813.4210525000005,938.5526315000002],[845.8690315,914.4629344999998],[833.6230990000003,907.8358475],[847.9513360000001,900.1584185000002],[525.7172709999999,935.3736065000004],[525.7172709999999,906.9534470000004],[523.9985769999997,878.5949945000003]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"338.41267","left":"489.86671","width":"1116.80134","height":"773.65892","x":"489.86671","y":"338.41267"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_8\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_8_0\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_8_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_470.0000000000\\\",\\\"962.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_1\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_1_0\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_1_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_365.0000000000\\\",\\\"962.5000000000_365.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_0_0\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_0_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_350.0000000000\\\",\\\"977.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_0\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_0_4\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_0_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1082.5000000000_350.0000000000\\\",\\\"1247.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_8\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_8_1\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_7_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_470.0000000000\\\",\\\"1142.5000000000_455.0000000000\\\",\\\"977.5000000000_455.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_23\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_23_0\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_23_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_695.0000000000\\\",\\\"962.5000000000_695.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_22\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_22_0\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_22_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_680.0000000000\\\",\\\"977.5000000000_680.0000000000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_12\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_21\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_12_3\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_21_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1172.5000000000_530.0000000000\\\",\\\"1172.5000000000_665.0000000000\\\",\\\"1082.5000000000_665.0000000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_3\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_14\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_3_1\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_14_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1037.5000000000_395.0000000000\\\",\\\"1037.5000000000_560.0000000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_6\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_13\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_6_2\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_13_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1052.5000000000_440.0000000000\\\",\\\"1052.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_4\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_12\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_4_0\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_12_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_410.0000000000\\\",\\\"1030.0000000000_410.0000000000\\\",\\\"1030.0000000000_530.0000000000\\\",\\\"1022.5000000000_530.0000000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_14\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_16\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_14_1\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_16_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_560.0000000000\\\",\\\"1142.5000000000_590.0000000000\\\",\\\"1082.5000000000_590.0000000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_13\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_20\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_13_2\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_20_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_545.0000000000\\\",\\\"1157.5000000000_650.0000000000\\\",\\\"1082.5000000000_650.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_11\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_11_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_22_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.5000000000_515.0000000000\\\",\\\"1187.5000000000_680.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_22\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_23\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_22_2\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_23_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_680.0000000000\\\",\\\"1157.5000000000_695.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_25\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_25_2\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_26_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1052.5000000000_725.0000000000\\\",\\\"1052.5000000000_740.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_26\",\"endPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_26\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_26_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_26_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1082.5000000000_740.0000000000\\\",\\\"1127.5000000000_740.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_27\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_27_0\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_27_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1127.5000000000_755.0000000000\\\",\\\"962.5000000000_755.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_1_28\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_1_28_2\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_28_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_770.0000000000\\\",\\\"1232.5000000000_770.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg\",\"rawStartPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_15_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1367.5000000000_575.0000000000\\\",\\\"1247.5000000000_575.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1\",\"endPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1\",\"rawStartPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1\",\"rawEndPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1367.5000000000_575.0000000000\\\",\\\"1315.0000000000_575.0000000000\\\",\\\"1315.0000000000_942.5000000000\\\",\\\"813.4210525000_942.5000000000\\\",\\\"813.4210525000_938.5526315000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1\",\"endPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1\",\"rawStartPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_1\",\"rawEndPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"813.4210525000_1073.5526315000\\\",\\\"813.4210525000_1077.5000000000\\\",\\\"1315.0000000000_1077.5000000000\\\",\\\"1315.0000000000_575.0000000000\\\",\\\"1367.5000000000_575.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos\",\"rawStartPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_1_14_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1367.5000000000_560.0000000000\\\",\\\"1232.5000000000_560.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0\",\"endPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0\",\"rawStartPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0\",\"rawEndPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1367.5000000000_560.0000000000\\\",\\\"1292.5000000000_560.0000000000\\\",\\\"1292.5000000000_875.0000000000\\\",\\\"812.5000000000_875.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0\",\"endPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0\",\"rawStartPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_0\",\"rawEndPinId\":\"pin-type-component_a4250f4b-b7c3-4cd8-ad73-f9c1a5eeffc9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_1010.0000000000\\\",\\\"1292.5000000000_1010.0000000000\\\",\\\"1292.5000000000_560.0000000000\\\",\\\"1367.5000000000_560.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos\",\"rawStartPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_3\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"833.6230990000_907.8358475000\\\",\\\"962.5000000000_907.8358475000\\\",\\\"962.5000000000_785.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos\",\"rawStartPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_3\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"833.6230990000_1042.8358475000\\\",\\\"962.5000000000_1042.8358475000\\\",\\\"962.5000000000_785.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg\",\"rawStartPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_4\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"847.9513360000_900.1584185000\\\",\\\"977.5000000000_900.1584185000\\\",\\\"977.5000000000_785.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4\",\"endPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg\",\"rawStartPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_4\",\"rawEndPinId\":\"pin-type-power-rail_a818362a-9609-419e-afdb-0484a3ad4904_0_29_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"847.9513360000_1035.1584185000\\\",\\\"977.5000000000_1035.1584185000\\\",\\\"977.5000000000_785.0000000000\\\"]}\"}","{\"color\":\"#FFA6FE\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_9\",\"endPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_9_0\",\"rawEndPinId\":\"pin-type-component_e856bf6f-239f-495d-9f01-2780e496b019_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_485.0000000000\\\",\\\"887.5000000000_485.0000000000\\\",\\\"887.5000000000_914.4629345000\\\",\\\"845.8690315000_914.4629345000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-breadboard_a818362a-9609-419e-afdb-0484a3ad4904_0_10\",\"endPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a818362a-9609-419e-afdb-0484a3ad4904_0_10_0\",\"rawEndPinId\":\"pin-type-component_846761e3-79a5-45ce-9f89-d8258e1f2e70_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_500.0000000000\\\",\\\"902.5000000000_500.0000000000\\\",\\\"902.5000000000_1049.4629345000\\\",\\\"845.8690315000_1049.4629345000\\\"]}\"}"],"projectDescription":""}PK
     ��/Z               jsons/PK
     ��/ZA���/  �/     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"2000mAh Battery","category":["User Defined"],"id":"2f403b15-90c3-4075-86a3-7ea6b108dda1","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"d20a931f-9d34-4029-b213-4c0e689ce6a6.png","iconPic":"cd711d72-4439-4fb4-bf4b-39cbaf4dbd75.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"12.32128","numDisplayRows":"16.29902","pins":[{"uniquePinIdString":"0","positionMil":"655.28070,1527.78699","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"555.28070,1527.78699","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"APC220","category":["User Defined"],"id":"cc6ddea1-99fb-411d-bfec-02f29cfc7b20","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"4ae07c11-480c-44ae-b2c6-f8186e930d96.png","iconPic":"fbc1041b-f35a-4c82-8c92-5608856c8a22.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"16.68849","numDisplayRows":"7.66768","pins":[{"uniquePinIdString":"0","positionMil":"76.08892,689.51916","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"76.08892,589.51916","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"76.08892,489.51916","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"3","positionMil":"76.08892,389.51916","isAnchorPin":false,"label":"RXD"},{"uniquePinIdString":"4","positionMil":"76.08892,289.51916","isAnchorPin":false,"label":"TXD"},{"uniquePinIdString":"5","positionMil":"76.08892,189.51916","isAnchorPin":false,"label":"AUX"},{"uniquePinIdString":"6","positionMil":"76.08892,89.51916","isAnchorPin":false,"label":"SET"}],"pinType":"wired"},"properties":[]},{"subtypeName":"MPU6050 Accelerometer + Gyroscope (Wokwi Compatible)","category":["User Defined"],"id":"70f88287-3db7-454f-a714-3fcb737f1bfe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"42ade947-84bd-4266-8f8d-47ba602ec33e.png","iconPic":"ec55ee1b-9bfc-4adc-bb90-2198f3917cd5.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"8.51653","numDisplayRows":"6.34167","pins":[{"uniquePinIdString":"0","positionMil":"76.35354,574.02468","isAnchorPin":true,"label":"INT"},{"uniquePinIdString":"1","positionMil":"176.35354,574.02468","isAnchorPin":false,"label":"AD0"},{"uniquePinIdString":"2","positionMil":"276.35354,574.02468","isAnchorPin":false,"label":"XCL"},{"uniquePinIdString":"3","positionMil":"376.35354,574.02468","isAnchorPin":false,"label":"XDA"},{"uniquePinIdString":"4","positionMil":"476.35354,574.02468","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"5","positionMil":"576.35354,574.02468","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"6","positionMil":"676.35354,574.02468","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"776.35354,574.02468","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LM317 Voltage Regulator","category":["Power"],"userDefined":true,"id":"0a0aa907-9846-42ff-9576-36638174fe13","subtypeDescription":"","subtypePic":"fae5eb44-bbe2-4b21-a13f-fb7a66868d1d.png","iconPic":"aaaf988e-4d8d-46a5-ae55-a0506af48a51.png","pinInfo":{"numDisplayCols":"3.69980","numDisplayRows":"6.23170","pins":[{"uniquePinIdString":"0","startPositionMil":"90.01000,0.00000","endPositionMil":"90.01000,-100.00000","isAnchorPin":true,"label":"Adj"},{"uniquePinIdString":"1","startPositionMil":"189.99000,0.00000","endPositionMil":"189.99000,-100.00000","isAnchorPin":false,"label":"V_out"},{"uniquePinIdString":"2","startPositionMil":"289.97000,0.00000","endPositionMil":"289.97000,-100.00000","isAnchorPin":false,"label":"V_in"}],"pinType":"movable"},"properties":[{"type":"string","name":"Type","value":"LM317","unit":"","showOnComp":true,"userVisible":true,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"SN74HC86N","category":["User Defined"],"id":"7799e1c0-2491-44a2-a64d-b6a1e1bb7939","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"e8fbe2d9-26e0-4ccf-9f9e-bb43371c63c2.png","iconPic":"95d79837-2dff-4c75-b12d-e13dc3081ed5.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.86081","numDisplayRows":"8.64605","pins":[{"uniquePinIdString":"0","positionMil":"42.77929,729.96514","isAnchorPin":true,"label":"1A"},{"uniquePinIdString":"1","positionMil":"42.77929,629.96514","isAnchorPin":false,"label":"1B"},{"uniquePinIdString":"2","positionMil":"42.77929,529.96514","isAnchorPin":false,"label":"1Y"},{"uniquePinIdString":"3","positionMil":"42.77929,429.96514","isAnchorPin":false,"label":"2A"},{"uniquePinIdString":"4","positionMil":"42.77929,329.96514","isAnchorPin":false,"label":"2B"},{"uniquePinIdString":"5","positionMil":"42.77929,229.96514","isAnchorPin":false,"label":"2Y"},{"uniquePinIdString":"6","positionMil":"42.77929,129.96514","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"342.77929,129.96514","isAnchorPin":false,"label":"3Y"},{"uniquePinIdString":"8","positionMil":"342.77929,229.96514","isAnchorPin":false,"label":"3A"},{"uniquePinIdString":"9","positionMil":"342.77929,329.96514","isAnchorPin":false,"label":"3B"},{"uniquePinIdString":"10","positionMil":"342.77929,429.96514","isAnchorPin":false,"label":"4Y"},{"uniquePinIdString":"11","positionMil":"342.77929,529.96514","isAnchorPin":false,"label":"4A"},{"uniquePinIdString":"12","positionMil":"342.77929,629.96514","isAnchorPin":false,"label":"4B"},{"uniquePinIdString":"13","positionMil":"342.77929,729.96514","isAnchorPin":false,"label":"Vcc"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Electronic Speed Controller(ESC)","category":["User Defined"],"id":"e60aba2b-e9b2-4ddc-8d1b-286ba98ca1ae","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bce349f0-9fdd-490b-ade4-f6d95f909232.png","iconPic":"4fd5fc97-bc4f-4740-9bc3-7af0136a9299.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"24.25450","numDisplayRows":"7.48979","pins":[{"uniquePinIdString":"0","positionMil":"341.22807,135.16840","isAnchorPin":true,"label":"Battery VCC"},{"uniquePinIdString":"1","positionMil":"335.08772,558.85261","isAnchorPin":false,"label":"Battery GND"},{"uniquePinIdString":"2","positionMil":"118.76786,398.25463","isAnchorPin":false,"label":"Signal"},{"uniquePinIdString":"3","positionMil":"200.40741,354.07405","isAnchorPin":false,"label":"5v out"},{"uniquePinIdString":"4","positionMil":"104.88583,302.89119","isAnchorPin":false,"label":"GND out"},{"uniquePinIdString":"5","positionMil":"2253.11293,537.65911","isAnchorPin":false,"label":"M1"},{"uniquePinIdString":"6","positionMil":"2253.11293,348.19138","isAnchorPin":false,"label":"M2"},{"uniquePinIdString":"7","positionMil":"2264.57089,159.13503","isAnchorPin":false,"label":"M3"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Electronic Speed Controller(ESC)","category":["User Defined"],"id":"e60aba2b-e9b2-4ddc-8d1b-286ba98ca1ae","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bce349f0-9fdd-490b-ade4-f6d95f909232.png","iconPic":"4fd5fc97-bc4f-4740-9bc3-7af0136a9299.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"24.25450","numDisplayRows":"7.48979","pins":[{"uniquePinIdString":"0","positionMil":"341.22807,135.16840","isAnchorPin":true,"label":"Battery VCC"},{"uniquePinIdString":"1","positionMil":"335.08772,558.85261","isAnchorPin":false,"label":"Battery GND"},{"uniquePinIdString":"2","positionMil":"118.76786,398.25463","isAnchorPin":false,"label":"Signal"},{"uniquePinIdString":"3","positionMil":"200.40741,354.07405","isAnchorPin":false,"label":"5v out"},{"uniquePinIdString":"4","positionMil":"104.88583,302.89119","isAnchorPin":false,"label":"GND out"},{"uniquePinIdString":"5","positionMil":"2253.11293,537.65911","isAnchorPin":false,"label":"M1"},{"uniquePinIdString":"6","positionMil":"2253.11293,348.19138","isAnchorPin":false,"label":"M2"},{"uniquePinIdString":"7","positionMil":"2264.57089,159.13503","isAnchorPin":false,"label":"M3"}],"pinType":"wired"},"properties":[]}]}PK
     ��/Z               images/PK
     ��/Z�ȅNܶ ܶ /   images/d20a931f-9d34-4029-b213-4c0e689ce6a6.png�PNG

   IHDR  }  �   �=:   gAMA  ���a  
IiCCPsRGB IEC61966-2.1  H��SwX��>��eVB��l� "#��Y�� a�@Ņ�
V�HUĂ�
H���(�gA��Z�U\8�ܧ�}z�����������y��&��j 9R�<:��OH�ɽ�H� ���g�  �yx~t�?��o  p�.$�����P&W  � �"��R �.T� � �S�d
 �  ly|B" � ��I> ة�� آ� � �(G$@� `U�R,�� ��@".���Y�2G�� v�X�@` ��B,�  8 C� L�0ҿ�_p��H �˕͗K�3���w����!��l�Ba)f	�"���#H�L�  ����8?������f�l��Ţ�k�o">!����� N���_���p��u�k�[ �V h��]3�	�Z
�z��y8�@��P�<
�%b��0�>�3�o��~��@��z� q�@������qanv�R���B1n��#�ǅ��)��4�\,��X��P"M�y�R�D!ɕ��2���	�w ��O�N���l�~��X�v @~�-�� g42y�  ����@+ ͗��  ��\��L�  D��*�A�������aD@$�<B�
��AT�:��������18��\��p`����	A�a!:�b��"���"aH4��� �Q"��r��Bj�]H#�-r9�\@���� 2����G1���Q�u@���Ơs�t4]���k��=�����K�ut }��c��1f��a\��E`�X&�c�X5V�5cX7v��a�$���^��l���GXLXC�%�#��W	��1�'"��O�%z��xb:��XF�&�!!�%^'_�H$ɒ�N
!%�2IIkH�H-�S�>�i�L&�m������ �����O�����:ň�L	�$R��J5e?���2B���Qͩ����:�ZIm�vP/S��4u�%͛Cˤ-��Кigi�h/�t�	݃E�З�k�����w���Hb(k{��/�L�ӗ��T0�2�g��oUX*�*|���:�V�~��TUsU?�y�T�U�^V}�FU�P�	��թU��6��RwR�P�Q_��_���c���F��H�Tc���!�2e�XB�rV�,k�Mb[���Lv�v/{LSCs�f�f�f��q�Ʊ��9ٜJ�!��{--?-��j�f�~�7�zھ�b�r�����up�@�,��:m:�u	�6�Q����u��>�c�y�	������G�m��������7046�l18c�̐c�k�i������h���h��I�'�&�g�5x>f�ob�4�e�k<abi2ۤĤ��)͔k�f�Ѵ�t���,ܬج��9՜k�a�ټ�����E��J�6�ǖږ|��M����V>VyV�V׬I�\�,�m�WlPW��:�˶�����v�m���)�)�Sn�1���
���9�a�%�m����;t;|rtu�vlp���4éĩ��Wgg�s��5�K���v�Sm���n�z˕��ҵ������ܭ�m���=�}��M.��]�=�A���X�q�㝧�����/^v^Y^��O��&��0m���[��{`:>=e���>�>�z�����"�=�#~�~�~���;�������y��N`������k��5��/>B	Yr�o���c3�g,����Z�0�&L�����~o��L�̶��Gl��i��})*2�.�Q�Stqt�,֬�Y�g��񏩌�;�j�rvg�jlRlc웸�����x��E�t$	�����=��s�l�3��T�tc��ܢ����˞w<Y5Y�|8����?� BP/O�nM򄛅OE����Q���J<��V��8�;}C�h�OFu�3	OR+y���#�MVD�ެ��q�-9�����Ri��+�0�(�Of++��y�m������#�s��l�Lѣ�R�PL/�+x[[x�H�HZ�3�f���#�|���P���ظxY��"�E�#�Sw.1]R�dxi��}�h˲��P�XRU�jy��R�ҥ�C+�W4�����n��Z�ca�dU�j��[V*�_�p�����F���WN_�|�ym���J����H��n��Y��J�jA�І����_mJ�t�zj��ʹ���5a5�[̶���6��z�]�V������&�ֿ�w{��;��켵+xWk�E}�n��ݏb���~ݸGwOŞ�{�{�E��jtolܯ���	mR6�H:p囀oڛ�w�pZ*�A��'ߦ|{�P������ߙ���Hy+�:�u�-�m�=���茣�^G���~�1�cu�5�W���(=��䂓�d���N?=ԙ�y�L��k]Q]�gCϞ?t�L�_�����]�p�"�b�%�K�=�=G~p��H�[o�e���W<�t�M�;����j��s���.]�y�����n&��%���v��w
�L�]z�x�����������e�m��`�`��Y�	�����Ӈ��G�G�#F#�����dΓ᧲���~V�y�s������K�X�����Ͽ�y��r﫩�:�#���y=�����}���ǽ�(�@�P���cǧ�O�>�|��/����-G8�    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   	pHYs  .#  .#x�?v ��IDATx���y�nYzއ�ְ�o:�cM�Ʈ�f�VSlJ�D��8v#r"	� H��� �����A`'�� B`
�-ؔ)Q�	Y���94�=U]㭪;�{��{\S�X��{�I!��,1�]�Ź���o{����}��}�!�d<OƓ�d��1�?�x2��'��x2��'A��x2��'㟣�$�?OƓ�d�s4�?�x2���_�����٨�DÍ�e%��p��&H�"��C�������N����~�'D��d���w~�_ޝ���Խfq��y��lB:c�Eo6��>����qe!�K�J��c�B�1JL�L�$�R�H2D�q���?ނ�d<��x���'���w�Oڟ��O�Ճ�BH~^$/-���N�M�v�0*)Y��2��o�%gd9h��&hq�D�L~��ɲ��P�M��m0H�%� �k� /��p2~��H2 EJ	��)�HF�u2��P� @��"� �r	����}�3l���م2>���y2���/�?�?����~�Ә��x	�I3s�C�	���d�m�ݗ�ۖ�dB��H3Hb����C?��L�h%�\k���XR��Q��$1���o�k�����2�2��Y�>wS���5!H<BF@��p^"��!�Y���g���$ɐ�9-rD!�Dɒ�_���T!��ǓL��x2~�a��u!k��k?����� @�� B�K�%]k�W����GL�a��C��|�Zu�l�aRI� Y�������o��;��"�D�
x�2�i����sD����!�B!����?1V{�	!������C@ E�R
)
B8�Z��s|h�2."&�+�쒧��uR�����R \9��{-����_~��)�'����d<6������ʋYx��i���B�=1�<� x]�P�-���,������<W$�O����C���=�*r�9<<��D���R|�� 8��1(�!|�>�8!\, ���_�c�����/�.�C<' �Ź)%I�`]���*I�IN�o�mJ۶�n�C�ǿw�v<�!������9Bh��Q�8;��`���O*��8>R��|��վG)π��+B`�{t�2�¯|�&u��o��R(E#�r�H���]�F��5�Z\�	�����f�7�B��`���
�<dFS��>�4O �[]��;���o���?x�pg/�E�W��Ta��@����!D��J@)J%x��:�19�hh�-���!�~���u�$A��@K�� �N"ZOj����[,>�e���)ӌ`/����APfxtN�e���!S°�/i���8 ��6B�pT�2��)H	 ZB��H=W��os�J�*C$�6��U|�b�O�%`q�=�s$���!K��Ւ9_��]~�W���5�;��)%�0#�9H�R�4MB UB�e�bU�RJ�p�INZk4�ӯ������_����tK���'��SE��2}�=��H�b�;�\J��K������,�Ya��T��R�*CR��m[�����ZKo{�tD���3�tTAP�.̑R��ɼ :h�X,T�$C�*UB�
�*TrN���uJ�p��!����K��!E�A�Rj�Dȱ8i.�#����B����Y�t��v|<~R�ӂɭ?��\|��[�Z�h��'��4N�_Ku{���s�,N������S��mI�e^ 3Y@hR���=H�Wb��()�"��Qy��"o�� K�1��z�21y�! �@k��G�Ĭ�3.2�G�C��'m����*�<
���qx���Bx�K�����=2HSҴ�cm���.�����9G�L+z�hM����}	c��{���4�U����<^���&KK�,BNB��,��#Bx�"c����-�*.�>}�W�bM�(|�Ǟ������B|�!�8rD(@��u���R�E)�L���?����HA�PKr5��!�Cp5"x��ar�Pc�-B;�B�wkr�@���Sh4P0������#��Ef����`�W-I��t
��@�@��Mx�>����n�|�I%�U�<<��N���:��뗫~,3���>.�^`�C���ˇTlfX�B��{ZӲ�,��x�ژ�� �2l�T"QY��ftV��)Z�Q�!�(�Ι����Y��L����M���g��'J��X��_N���v��;/t�w?[m�on%�qxmy���	�H`���&���A�nB�Z���! �"�+!�$ =/b��d=VJ��9H?Aye
��4І0�S|�H�1ɰ�қ��������>؀�6h[<
�H���
��# VE���|�"�Ü��j@}�b�m\̂��kX$�G��=Z0� ���N��*Tf!���m"���t|��D��J<J)z��U�UH'����s��{ayP��lɲ�nZD���ӊ=A
�뀠2��!�Ż$VeA����	��5Az�L2@ѵG�%����ދ��P9)��X\`�v�Ib�(R�)���;�j�������&��L �k���K�DA�u�yN0>x�8��Q�`m̆��:�5m\a)bn-D�5���ʥ�1kh{\�B���ihۖ4�Xk�r6����K�|Ӣ���sK��$J�!��Y|���8n��!�s�T��q8D��UUQ��eCp��Wv��\LB �=�o	��T(�"X#�Pn�+���ߏAF臌�(�d��gշ�g?K����#�J�����fR������y��C_���99ya]�%O�@��^p�V��Ա�T�;o�t=�pr!��+�II�8��8)��cЏ��eFb������4	�4#+=���{?�&�u�l�d�;��@�u��J��A�,�_���?���[LD �p��L6���l���8�G�| ��ه����?2K��{���W�!�`!! x7���	�R��"�:�	"�x��Wo���X������f��z�l(�B�4aH���k,0&�2t�)˒lT�ZOe���0}Go|$�u�w��Vx� UJ��H�G�1)��c�A��4Y��e��iX.;�4�ǂ���*".8b@	.�q����4ϩ7��~���������HA_:��M�=:A>���g:��@�,��`+`�m���w	);d���vC��%=�	���&D,k	��V�؄�VT�@�+���;l��"��;��&)�.�6���<Z�B��Ah0�.�!I.2��"�.R��TG��R�	�6�Q΢Z����q.0R+JA��!C�]�A�/,"�ٞ�c%�6t�q� <Bx��6dY��EPY�T	���JTVDN2����ӧ	">�R���n���˧��>�ډ���gH������̟����ܿ��x�w^6�=��W�i��p�uk2��;�v�O<��+���i�[׹��`�3����?|NN�g3�{r]�>�3/!K@�(�b�b2���I���P!�ڝ����|p�|��矇g�j�&(��H%I�A���wX�~�t�2*R9��kL���ꋠ��Ayȗ�4�|��/��0o%v�F/~��x��� ?�x<�@�1���7��0��=�ޡ���#��O�e=����um��4}o�E��ڎ�+�\� +=���B�$�S��&_R�Y�C��W�I� H�a\Ke=Uա��Ȅ"��#��b�H�*K���x|�2RxE3���S�OHC��!��FJ�
���G(�k��H�"d	!!�-�ڥpJoa����~�_�g�?ZЗr��yd�ưl�l\O�kH���=ֵh[�\.��+\X��b�a:��� ���%$=B���'��644*Є�5���$.j���e��rc�y�t:�(�Ղ>@Y����\?3�%�i� ���F#���V+�2 �RBlmm�g��>m�"��C�>�S9Bq!��)
A:,(�	��H�RҐ��Ib&4��1�Z��ò��9*+�ɘ�Ag$A�$�!��;��H��<�w]�Y���!�N�j�����gG�"U���^�{�>�y��wb����+b�&4�n},Vw�9]�~�|y��e�wVU�J���;�.VdM�'nNp��:Ǣ�4��`�ܰ^KR��"�(�6k����d�Є�}�w�@�H&�	�uH�o'<NB&B�2Ĺ��AY�	R���`�^D����O�}����}޽�?���)���~v��
�u�^P�N8;z����kۚͦkb���Bכ�F����9En*^_).p��> Dx�����G/��E�|��P'\�A�!/�Ԃ%IR�E�B
��U�1�����?p}���#I�U�՜ym���:p%,[XwY��L?\b.�g	:�/�wk.x��HҜ$�9�{��$MJ�d��:�Ν#�f���4T,�!R8�n�j���#hAi���G�*��IB��!I�W�S����A�ȇ��&�����������ӳ�@,�9�4�Y��u�ċ��i� ��H�Aߡg��093��c;"q%-������X�q�n���U�(�]���`>^Ҙ�r	#;��W��I�5�\��l������[��]�t�$=AI�d\���s6kOgJj��A*�B!Z�7�p��V�Of<��)��� <�№Z`Ĕͦ$ta�L(�1����*�b�$͡���5� �M�J�1��"1֤-Y�V�h�x��rk���c�lɦO�Z��6!q�����K��!�d(��[pz�֚�O�b=��+\�A�����8D�/�Ë3���r���f�R
�V�����'Ha����Jd��}~�M�?x�M�p܀
�Y)�6Ι�K���~:�e��zM�u��hm��
�����㾽K�Yv�
O�'w��W���+�i�[EbW�>���F7TZ��rH p�,R��!f�/!	�X�$����\h����_��۸y�l2A�6�9�6��	!�"�D`1�G�Gٺ �,b._烸T�Q���1r��E�ƤdVH)9φ��92$IH!�UT��a�^'�ٶ!
$4J�s�x,(� �E�%B
"[a�4�L6`��ʀE��)L"�9]�pzz���z�@���QB�Ņ˹HZg)��!IL��%X"���P1)I�I��tȐC�Y��fÝ�E��՛%��PN���m-�U�T�8�%S\�H��H�9e~�:�a������F��T��k�;��sp�À�8�s�-P*�k���m��#/
)蛶E�>8�s�}���<�Q��I�ږ��K0<+~��̣ﺘ��8�T�	�B��;N��tH)�K����).IW��Z6��Ś�����P׎�Y�<��c8Y�0�Ab
֫��4!I�5�<EQЙc�%Q�\`�� L?x1��ӟ�V��F�)-''�l6�%�r�$(5pb@K�|g�rc�Nہ3�x;`�ֆA�a�E����Ef��dYFۂs^*���@=Zfl6T"HRAUE�V5�Ȥ�W��u(�DUo���z_�5��U����d���������	EQ`��w�V�8�h��#Kr��Z��{vږ�[�e`c,�����4�:qhg	�� c�P������1����޳5JQ�!����[��3���m���8���5��a�C.RF|@��_6A]H#]�Bᠮ988��w��4���Y=���Q��I�R�Cu�}���((��]�P=}Hy�(�\��s~��=!Z���хH���z�u3 ~���F��[w��UL�0)s�k� �"�RF#K��{�!K���SK����5��+֫���̶f8ב�e��B�Ĉ��Ϥt@I�*�����9�ȡ���}��sΑ�)8�rQ�0,���GG+�n���S�Fշ3�p�2�D��P�(�*���D>b�������92M�s:HҎ<��b�~�Ƙ�\&6��~���')�o��D����;K��b|��:BxH&A	�i��M����b\�BW"�h��H�:ÃUGc��O��](p�!��Q*E�G��+O��9�)9o�q�wy���nx�+����k��7�>�4[F���<��2A�E�
����ヮ5��F�d��u�>��6�i��=�Y,a6S\��c\��	]�x.���)�(�Y`M�t�u�=�Z�$B��s��fc����,��<�;_q?�D��ڱ�A*���p��W�C�y��D�\gAKB>CxO��H?P5��~���3\X��)r��R,Q���x[�����C��(�q�͢���iiQ�"�2FuK�wt�9�W[r�iC�hi�م�_H���824kP&���w�T�b�s����=���-�>�I�DA�=����Y�pS����=��d�0�Ue �@gRD�N\�c �-b��{���;�����'<<��h6�F��J��)�ƪ���x)�*f�Q�#�j��~�R�y���V�G�q.�e��/�Ђ�m�r�p�V��ݠ�o�IhUL60��r��;�t�e�R�H��0aP��1m��N��l����X��c�>e>��W���[�X�ֱ;B
��䜠u|Ul�� �^\H�F����-�H�j�1=��ɍ�4��a��(�	����^o9��x���c��CFɂ��Wg�BZ`��S5A���S��"�8�G�w0�w�"���	��$6'ȇ(;���H��	�&�@?|������e���G'��)t�v��q1�?��:*z��$IB���ީ�����=�͜岧J0����%!��b�bi�b�ӷ9�eI�$x�r~Z,��7���3�}�c�6z�L*LlmD�t�u4�����5y1�$�x�cEY�������9=��i�YY��x�cT�g����p�j�d�Ħ	�IMH�(�0���NbQ��Y��}����q e`�T����h;�=���G����f�L:���k�����nI�C��p���s7��U��YL��o��}l��+��.Ù��h�l��$(���=M���}ݬVL�StU�4+�IM.�����r͵��+{�IG��^
�T�C9�Z�t<��[[��l��-m�	FҺ���B+�
�д��K �r�2�-ݦ&���0��4Jx@��Cʈ�{P~	<�YNNN"f�MߠT����������)�%��A� �� �#9��Gā���B�~��vi��9��c���(��C�z����I�A�de�j�Vx)�%Bx��5�"PhKQX�T�c��4x �_st��^sT>�E��Й��]}�.��gR����t�%�Au'�u�:��m�:xU8��Kc:�Ҵ�+�ַ��r���\KbO��Hi#�%<A���{+��"����'��˨ܒ$dI�H12(�R�a[C��H����?z|��߄����'����W�mld�Z�Uw��Q��v���$Y�!'x�i�-m����sTI`e,��t[��P)�����A�s��4*�����i������t��OM�̮if/�Xf��ΘnAVXF�mN��YPZ⽠kM��[��
!=BG���Бt	A�e:�0;�Zsz��^���t����JJ���;��b{[1.5���<K�����d�\4$�'�(4�'�9��4�S�8�u��Qh�b���Vx�X���4�������-T�Ԇ4Mu�ā��TEl��70%��T���:C�)#1���yʩ�����clGnj��u���t�Y����Y8I'�z���6Xux�t�넑8��7�Մ��H28�ʒo�����c�;���L�x�ݣ%��;�v�!�V��Yy�%�w�D;V9������A�QD��@���j(3�7��9z'�2��Qz�|4ES�N^k�f�����9�����:D!��բ�$u�0v�`� P����� 4�1���	�������!�b!�"F�>���5�}<��� fXh�������ItJ�d8+�.M�ё���,�ʂ���5��b,˄;���x������	�YA:�c�bqV�G&r�c�6�����،�A=\)c�猽�n�0��=+&s���L�՜����.�h3''�Ta���k��
�i�R���G�44Y+F�Cr�U(S�oc���BC��|4"�w@vm�=�a�nՍE��%\_����RgR9�Z\ߡCl&�lċW�9��I�E�14M��b�mGG��ԧ���E��:�KX�V�}O�u�a;�3U��H�)�ᔊǩk<x y��aT�<�����m����o���~�:g'-˳s�}�/�_���9����JH�4v������m���:�߁��z� �g���X��ް\�l60� �����{�;l�P��/U�"#�v:c��x��K!a���1�ٽX�
��b�`{;#$�hZ�Kd�І�k�
rb�4T�h��3l(��#r[RSI�K�(�G)A�6��5����U����X�%���M��>�X�5��u�S�5[��7�R/G9Ũ��c,Z�l��@$�����)')��4�226�HN�����
�H^_V�n��*`6��q����&�R��r� }x����s��H1��ȣ�#��a�Q3=���x�)�����?1�+{���(�3�р��2��U�~1�ނ��`P�X���*2��Ts��K���Z�-�H��Ӷ��E@�!#7a�QB��l�e��z͢ސf�� DOm�1����I�BF�K���R��	�Az-U|^�p���R�&��}��̢��{Db�sR%�����@Q$��,6Xt���d�(�v.> ��И�m5��%�@8��{P	}۲^�Qml�������q�$�#}�<��}LA�dp@�ޕ�VdE�r�`%�{�Y��n��=ipI,u���'q�D�tN�U�[�l���Rc= 3��:!ͮSUg�<6�=�"��c�����2���v�?�E�s��g�_P[GH��[�6 !���Xbi:�cy�T oʢ�kc_��o�*B'(�uI�j@�U����ЇQn#�)Bz߲I%W�;������6p�{0����*�Ns&[� �IӅH�;(&P6���d��<蓎�mgB'��EvqR�CVkᚻ1�wǑ�k�kM�G�r.ֺ�oh�CG��e�y^��a��Zh��ܺF۶L�s�L���NsN�|I�5�z�����s3DWѭ�t�S���w-�臐�y�Nѫ�W�#|�u�Σ{�j�	ڂ�LHa���x�r��X��;�|���rX���޴�"�Z��R!��'`C��
��:ҥco�^�����Ë�^+�1��G)�����d��D���}@_$Y��%K{� A�C6�[V;rK��*/c`��4�1�b�o�(m�$��\BzA�j�Bbd�מN4FZ����fG�F}~����!�'kd!�ik��d���@�H�n,��@ I�%�om�0����k�q@M��F=��/ZP�8��n���.�Ś�jq�%H�ښ����]���	�\��	��|�s�o���I�DȎ �N���..�M��>:��*�h�0r�{�^R�1����/�G
�Z룦i�KE��D+��13��lD_n�&HJD��C]�$ސd��Hqv樏����H�{�!�ݴmlm��°ː!�9����\k�������h���c-�ǂ<ϑ�����K�˚ �F)K����b�ԕ��<ϱ}dߵ�131QA`6�Rlo�r��l(vc`,
�IBU]E��ɕ+�!�ڞ��s��T�'����E&1ؿ��7o��l���w�g���s�Aˋ/^�J6�?|����7$tdY�6�ԫ[\�v��Ն�~�]>Xh�\��tk���9���MGOݸ�+W�pzz���=d�Z1E	gSEl>�MӰ��H�4v%�;
׮��,g�)6RGu�����P��8集j��~C�h@�3���x>�����xfBr�:�[oP�4�;��S��}>����Ch���'�ne��q `���r�m��g*��'8�d��ݦC���km�|tkY�!hR��(8h*Z%H�Fb�/b0s6���ʫ��]��p>Z�x�ڋ��G
1�JEl=�K��e��^�t���8�=@�Qm��^�߿�H���ݐ���H���p?y%dY�>�:\@י��iy���ј����(���1�%�N�����m��a͵�1�bA�i�V��#���{�(-����$IB��D�.�Z8�x�t�#�'�K���]�	��hDȹv�)���9��Grh�$y��m�rE�$m��,�P:���V�~�"]dY�P cX,��>�r���E��X65�HA����������SW�xk�Z�� E�YF"��X� ��g���e��AYAR����_6�E�=�(�Z�f�iz����G%��@B��
��}�7�Քg�úo�jp
�ц�x>���:�Y��)L�n�`�&p�ʄ�Ba6�Q���MEJ�$6��o'Ȥ"��4���3�h��*HB�
�SY:C�R���o���\o,W��H�:�pg��y��
���9z�Л5����t�?8nЕ�Om-��[��[-�>?���Gz�Eb,��7_���Wy�w�ҵ��O���n˕mǫ/'���7-%���t�������套^f4}�����ß~���͞���O�hv#n�4sv3I.=���t���_fkzƬ?��gs~��7,����/Q��e4N��+���߸͛�@�Z��t���x�S���G�o���Ը�y�u��܏��]��Kɢ14�)�ް7	L��S�
Af�Wӛ)>Y��)i�
��1�ʘ=)����,�*xo��ϥ����OE`��� x��Y��C��T0�B���	[8�BꞱ��<���BBQ�Y����r���G^��Q���/�X��Ï��Q��}��#�K)�t`ZHRŴ��3X T*.��
U���"���	�	A@UU�:A%tU�t���H�EJK=*�eOV�x�����U����&�+�&c���e��Jut�.]�$՗v�D;e���Jtppų15��3:8U)�t�ҁE����q,{*m�sƫ���*�nC�*�l_�=�mO�&�U=G�5_�=Z'4�S��X���L��64=dI�����H5�X��?�1ʲ�2�Td�75!2�������V�K����mI.W�U�#zO1їD����O����}�OU�!��Z�c���l�4��d�ã׮�3�<�{�o��;��� )�:�l�2���F�WnJ2(G����=$IM�&x����Z~~�����E�Qj,��� ��(���P�	*�}o����-�^}��S���loNO+B�F#�k0F[Q�qr2��"��S�v
899aw��$��e�X�V\�ܼy�_�;�ʷ���yf�d�����٬¹#F#�N�\��y㍚����q{;��e�E�t��x'eYB�x�|~��z�;8ӑ+��,{{����?���؅?�'IӔ���:vc��]�3��{v�)�k���*��� ooa��ԧK�^#�b#G�. �:���i��ͻ�(/ε��ɗ�Q}��{V�y?��.���� k;�QݥM>g1=�'��C�p*�eJ&�1M�{{����#�~��ͦbg4�0������^��C��MW�~����B��`/I���@/HR~hN8����Rn[(3��h���1=h![`�~�BǷCU�H� u��꺦G�$H�����q��t�����r�Z¥er �u@�3
5c-V4��Gk����z�j&QN���1q%HH���]�x"���݂�,�i ���x�v��(`2�j�ewVK�;�$i�jb<;�q��AW���,���<@e1OHR��gg8�8?�HUq-�KҾ,Knޜ����8'�s�M3�D���G�jk��yJ��Q��r���I}s�)$��_�2)���1:6\�)^	��1�JY.#ɳ<~�L�������{dg�Y���FB q9X��=��'��g=/�,����d9�+�o��ZF׭(K�x\RLUu��1�-�ygU�ۣ�Uw�1����f�l���,��ci��HRm�$(���Z2	I��`*P.p����sptN$�\�9�T<8�iV5���F�+k����P�SO/x��	�Æ�Y���ck>�y9�ڌ��#g�4�p2��m��ʆ?v>=>�F����g�
��˯q�}�d�/�Zq���>�e��_�T����^���?���i)xpv�Ͽ����9ree=|p����?�e����:�t�	c�{�U`����z½;R���dFR��g>u��T��|�/�$����s���p���#ʑ��6��.[��ĩ�S���999A��r���wVt�#I�8S\�z=�h��d�V�Y����#�h4"�$h:���17��:�m1	�$�Wom%8�!�F~(����#�#�=���wqɇ{D���� ��Sݳ	������k�T) I��E9 ��t³�=V��s.b�B�E�P��,���C���.��xL_o�-�rA���*�����=F��P�j��^E�©��ht�0��h9�+�C*E>rdY�R�jSG�'����f2�꠆{%���>ǩ-ڳ��9%��i����=Ayt��yK��l� 'jC�v��0yukL0ދ}9�wF�]�4��Ç\yƐޠy󵨔:x��
VE+V��MkVN*�:��-�t�#D�G�c��m�@�	xKp� �&�f �>IF���_�'����㊨a�ٰ\�܎n����w�9�J��1c���q��n~����%���W_���6����|^~y���,:DU�㜊D� ��L2�MTA�,Q�����97��X�X�Z�c�>r$�:��
�=v��7M�����4�R��sn`����m9:�[�rn޼�7��&�%��n�V|�;p��7�z/�������
���0�������>��S ��=g�����������{{2��|�C�&�/L���3�����w������}:#�k�n�y��~�N��m���{8�Dp������6�i��gg����k�{�`�������s����<�|����b솓3ϳק�}�&�*	���{���/��[O���%Fܿ���q||���X�/�l\�l9Qbgֽ'OrP�t��~-��gX~�������3)جE	Y�]���f�����w����������?�/�s��ip.G�G^8����q�Qx�u���T���<4Gq!�~g,uo��l ƃݭ��	ڦe��T���������1�cu�P�%�������m��������F)J%qG�Aa��l�bg���GNE��
8��%�e�R������{A�m�,�m���\��5_�h4�s��dL�u�f3�C63�9??�m[ʲ��*����t��F�Z�b�ڊ��vݣ=>���A_Ϟ���&w#��`�dP�\�ebg��)I�3�K�j�z��`m�A��yc�aD��ņ^EYa0������7��}�u5�wv�xz�i�p'��w	͈���߃0��_���x����7<�5�B����}�+G�*"1L'SV�yZ:F�y�b��!��|p԰�Θç$�QԽ�|A;�`��UF�����kB%m�
l_ ��Zrk˱�
Tȑ&�¢�	^H��췇��!a���W[~ꧾ�ӯ>ï}�;��k
&pW9� ;�i�A%�]�/>}�?{�P^��W��>��0+��;;O�w��Wx�A�(�@��I�j�7߅���s{��������=x��y�n�XgL��$	�rM�Op���эgd����������_<!k�{p�Y�xnWSH��LӔ�����mok�s�ʩ�g���L���O��ӎ�^����]R!SdVk�^�ܮ׼�/��

y*9_wt'9�VyJ��Y>�����iuB�����?����)<�l��VO�L��H}�0��я�A<�:e6�(���$QI%��WL1�$a��������i�N�qB��$�FBY
�$�`p"J{�����*x��)pa0���TR�*�:b�O�$:�4=}�˵�r��d O������-R�(_렲S��TU�fө%M%JG�f�������$x��'+$��u�<ѹ�����{rU t"��ϲ����L�i�s*[q�0�:��A�M㙨]V2s��]�j΢)�����nc�.�V��R*Mƒ��� ��6��j���zI�Q6|t2x�����p�||ǟ<�/1�v���F#ʲXr.�}�"�B�X�}�IB̄����3��/���}���.���0�s�2�?����.J)�2��驣i"�;t����W8�.;�ʲ���p��S�8<L�"899a���`��e�_��p-䥲(˲ة{�i�=��!vwglmm1�LbvB�(
��o|����b���|��'����7��KLP�x���f%�����ܻw��i��7�ɷ�}�֑3����
��~�
�<�o��zy��ש*X.���ۼ��}�2�F������<�e����U���;���㟞����{��?����'^��%��G��=eY^��.���hĭ[�b�*.�>�����g��١�{�z�&Z�b1���#6lo�l6%�����[o�f�^�4-�oW����sf3^I���t��$�e�Da�"6m6�![��tʗ���n�z��l6�MUy>��!SV��}�ĊY�:Q�"����瑋��=�ۋ��W�Lt��9����U�1�L�dx�B��t�������vYz�qn�e�����UU�[�qq��$�ڨ���N"a}��,���a�<��}Q-���)
M��X���Q��{&�	Z��EU���%9Z�������(
�*�c��N쪊A��CL��j�"�������eA��d�h6C�j����y�q ����"�Ap�FT8���c���岣�@�1i2ÚSl�E�Y��F��|���GL
����zB/i�k��Cn߾�Ke�Kζ�]A�B��QcPmK�s�N����/���Y�Q�uW�sm?�T��'�<��j1��-r�Ԉ�tLݝ�^�P�{�:�;���G4�Ck������/x�pJ�lQ�+�n�6�d�oh|��5R+�l��a=sy��9&£m`o{I�6,̄3�
&{S���n��,՜e�u����%<�Śt	�k}�?��G����AK�^S�1�J�{��
�(�+�<�?x��C�9�w��9�ۊ�?wd˚��S������VA54��c[�,乥�K�R�K�1Bf�*�s��U�y��krc���^EA]U�b���Ϟ��s�|���h�L+������{���쌷�lk��r�ާ��0� }��t�9W�综����|���i�#)5))������~f#�X�B0+6���Rq����n�q�~@�[v�yL&p���|��7�����E���J�<.굇T�Tx<^�Kh4�h�����8bp��)��*bx4�����3�O�,�U��Z�"c�7��8����Q�J4���̘��r�)��6!x��Q&�'-S��5��I��=nӠ�E<ǲ���[� ^Z�4# �o���~�	�Ӧ�g�#(�P���mV�bQt��Fz�E�i�J��{�>�C&[�tّGBO��5P$J(�K��S�-28z�RL� �Uƍ�-Vx���'�F���U� ;���퓊�;��v����y�h�1�\��X�tMͼL�i�M����O�OӔ<(t*����u�-�Kv���YZ�zVh-�NO������}�6\�:�޽{\������=�=v�/6i�C���y��q��R����~Ŵ��)z��3�2d/"f��sx%vP�u�ݝ;5���[x���t�s�kx�-x��]��4 7��-��Oq���(���Tt�$V2�2���,=J$`�C�e���2��*r��f<�5�C�gz�d�І��c�GuD�$,��ՃC������}�����4���r�d������H���4V���k����}�}�9x�����Ա�H���X��I��5�u���I�C`q˪�l6�4g�X ��Ν��]�~����f<�*�7o�d��;��o���s����u�x<f~�������#o��*Vr������Lk��sV�E6�!��,NN��!Im��6�R5H�z>|�spzXW��4eS�4�����L��7X,8�	ah��ͣ�9����b%��\?ڮ������֞���|q���=D����z�$����yt��ޢ��:��.ri��FtZ�� �"O���9O[�L&����ɺ�����Z�<Vu���3�FEZ������;pxą,5<��Evm/3��U+���j�؈�5�-G�z�k�:w��_T�q�-1���I��<��s�����ק�=���P/Z�>v�e�|�������e%e��L�(��2šJ���T�~�c	�]v�ļ��Z��ɔb���e����(��#q:v'��p���ۖ+W�R3_�����+;�oV�z������ק<\3��bBk�EK�<�{��"�`w/��ݟ� ]F���@+`�v���N���i�qI��4��	x�X"\��&�[o�K_��\�P�p��u��x@\�bU�V���%��I\*�o�H9G�	Mh�b���^M.T#N���4y�E�x�͚�o����-��g��$2F�%���u�l	[�����;��Ŋgfc�7��Zp|R�ҧ~��b��s�A>'z�Г���#����cm��Hk4���B��z ����7��#�&)m��dpL&�Z5F��s��Ɵ:(�������z���Nz@�=��_�>~��_{O���ʟ� ���h�������@��3m�^�����{oH�gWE�z���������)�s��c_Z�D��|Dc���K�tTp��󶃷&S���Wp��� p�6���[^zYr-�]���'��5���jk��+[|�\�k���O��l���F�K�T�΂�hU�ՠ��*�h��0>�4(��<�0�#ZM�EP2����Gp�T���L��u\����I�ӆ���?����5�~�����)"�F�Ȁ�>v�z���*�3W���xptΕ ��1N 8c`y:'�
�zjP�����[�Z�̱�c��$�eJ�4db�֚�]���+t:�[,Ť��kV+�L�	$f��p��`�f�e�\U���Σ�<�5uS3鯒�%s3G-zt.���ؽ��;'<��u��;T��)wm~DV2�a���O3������}t��@ڃ+p}��)��![zw7lĈz�kC��8�������BC߶-~�ԟN��K�{vww/1���B�~~�|>��/&�VT�|\a7Cj1�X�=��a��fb����x�w�nry��.\���"I��j�'�3��w�����`��,�۱	q���0�d��4�|�o`�ek�K�����n���0d�	M8;;�l�	!PU�<M�.Ƕm/�b��P⻁�T���Y�q��N�<�ܳ|��֭aË�mvvv���k~�W�B���s&^c�Q�E�8Or��Gb,��rY#�d4����7��|�s�b�Z�[�p?������<���
��c���-
.�Yy1���W,�PU-���0}�Ynܸ��)��?�c���������(���Ȱ��E�w�y�]�0����yN��1�,�.q�x�5�Q��Q�4������i����y3ck+V-B�4���.�e'��5\��q}Y�^`ձ+W����U^b�N�[u�_�@��2�qH���߃"rEQEVU\V/�e���op��5��-�o4���Ӽ��c��^x�s�=f��AY�ܼ��f����������̣������De�a�h9=5�à�[��4,q'��lI֎�����b������z����lZ��n����1z�u�J�Q|�C���(�B�Bau��߸q���; >�l� [�"����0������fC�u�<��36&kc;wt������?�O�?4>�L��#�%G?&��lv�r�i�d{R����iL�ê��ޭ9��1X���(��lE-��r�!���~ĕ�5��;lY��5d�.4;
�cv������c�`HҸ9H�0s	�\�o[ƹ�E�;|����ai�3���{��zLe�!D��v�d�̆���^qx8Bf=��9o�ʕ]D8>� �D'T�A�N�؜
�f�4��Ѓ�`�i'H� $�%���%�m�ʌ�mX��ɢ|`����<_~)p���_���i���w8���ٌO?�q�����?"�qJ
��
!�-���%�|$@9O(y^ ?�������/H��O{&�w����g��n#7�G���{MQX
=g��M:�`*R�0��w���Αdzn�мybQﭹ�V��N����<�ܘ/������b����УSC�i�2�*S4	�d#A��{|�ق���\�ZNO{�����{��1�+����Ā��p�dM1{��@�˜L�g%����8�=�����6�U�������x_��jS{��U�1����������K0��ǀ����2ZoG7�4�n.��]���ң�o-�J���ϥ�X�@���{�-8h�3�W�SC��٦�f�bρ<kȒ�S:���,�^��5��P;C� �j�\(Ί�ʷ�g����� u�����w�㜮QtCg��3�i#�&D��&�u���w	�m1���z��U�q�m(˒�6ԡ����Y��5.4�-��q]�q*���(�B�"�8�X���t��\qc�d~r��aw�9?�%��-��E��8���lz���,��
dHpA|���^�.�bV)'\���}��c��Պ��ʼ����v��1�������?8�j� 7,Vs���2�MY!ek�%%$e>h��~ӡT����=��Ʉ������ ���̴c<c�a�^�-cJ_x�\��ʉ��幆���$,u���hȾ i�rK�\�zvw3�c���7S�\�^�M�GJ��/��a��Dԧ8��U5t�J��Ƚ��!�$	�2f]M%�ؚ��x����o�x��C����_�P��d�!I����CRF^�ZG�FC�xL���9�2�P��=e{���Q�Z�]��4�=���_�|�g����ի���S7�L@-a�i��X�]d�u�����k�re�O��O�[����~�-�g���O��w��:a{{����z�η��h/<ib�7n����{�ǿï�6��g|�W�\!��,k���В$�����(��ei���=���ɭg�W$Ͽ�<h���}�۟���)��uk��8*�.��B\��v����UA���zi�&%Jz%Ȕ���C������c���~*��xꩧxu������s?��w�ܺU���ј/�J�<���>�R@obp���I:��t�����;䰷n��E��[>^��8����]H.
u�{����'~�Ѵ6ƋNbM $JI�|�6�Yy��� ggg$i U6��8�M�U��q�.8/�ݍ���F#NNNH��_4��l6���G���u�2u�ڳ,#E�q��E�H>�-@]��^(�.	{e���؂�p9�S%�4��7	r����U��o���5vnr6�E�)�:@�7�:��ă�S��)eN6*Y�9k1���sHy��t��[��ܸ�Z	V+�J@�
��iC�ؠ�6�UW�ӀD#M�v���RжTv�!� �ElK3E�4Y�f	vFP�s�`z�"������!��v�8o��ጳ%����[���	Mۡ�٤�l���L8>��^ԌF[�U�FiVm��4�Q*��IS���ӥ�>�G�!G�i��h���?���a[5lzIz ��
�9H��^���� ���C�G���1� ���$���t����]�݆�V�NRr�����}�N���'��Yx��@���]Z�v�UlP��؆&�<L|��������_���w�mS^�\ϗ>I�J�؆����L�ˈ��VF��i;��.�\q=���))��D��ls��6�>�[և��(H�ʳ��$�g0?��C�~��������~����c�����s>_�nHQ�CʞI�n���d��D"�YvCK��d�A���t�Q��%D�O�:fX4.�܋�2l�K*z���p�q�x�vK�^[�g眝���R��)���9�����Lư�JJR�b�T��2)@������ōN�D7�OUF�k��{hL����D�R�z�BÕ�G`3,b>�Q�S�C�\BwQ�
YV��г��Ք�F؞D�H�ɲi�*ڮ����� P@�������w�&O2F��� �YE���):xٲ�@��m��F'�2S925(Pz�%B'�$�"�ۉvMB�G�#hr�q��/�FQNq�G� ��3���G�v�J��#����b�ы�|<b�Gx%�q�E���f�{��ڨ�UJq1��{�=Ҧ�Z����Ƴ��?�,��#��ڴt�a2�P�y�gMq7��<��F$�DK(��c���"��,ˢch�P�5�A��1_�Zu��X��4�@ʻ�$�o۶8���f��}H�ؙLT�8��Z��{�.rE}N������(QQ����^����o?���όx�9I]ל�D�И�G�y�t����X�?d��|�ݐ9K��&v%�����5~o�I;���s���&��?w���8==�2��~���Y�sQSB�,�-����{jw���R�%x�J�(�ka{{���.B�\�H��[|gg�矪_݆�P��\�gw�!�%v-{wv"~�T|���pn�����ݚk;9�;�������˽{pm>�}6gs����O����~���h��>����ދ���r�+��T1���6�"����N��  ���k��^�b�����H ��a4�q����s0���.=�(
l�"��x�0.S|�_��1Hy�B삇���I���,�������%S����hAQh����@��'&r6뚦i88�$BҶ�`�NmI@)K��<.��,^�E>����iFߺ�s��wWr��=6��TQU�K�B>� _�T��(����B5x�ǁs8c�]��q���L_�HS e���6���$��h�3_?����z�b����{�:"MS&7�a{���	jT��̲�}
Jӹ@�Zj���Q��d���|�CN�?��7����+,sEoA����g���9-z0�f�(��~��j�đ�48g>��8�%�~�fcI�J=&X�Yv����b�f~z?�`�a���Ni��w��6i6%����q�Ԓʄg^�4�lϚ���������(!M����z���O�-�]�$����Lp�����v�Avȃ�cT�!��[3��*%�.6�dh��E�E�ر�W�*�(�H�b��]���1G�q�i��Y����|�E����xŝ^�=�G���(�C�uW�c�|e��/=��Y��'?k�ٟ�Ϲ�"�I
�i�6Op�����
�Z�����J�`�`�S;_^���E���Ã�?�?�$ُ;�|��q�����Q�B�Vu��會tһl=��y���G�y�5ig^}�����R�]��?h�p�5�2��c"� M2T�����z��CR3H;��m�C�5���@9i
��᫔�0�:~/�`1Xېs^��\��M��D{���w�s]�٫����y�wއ�Jh<d�%K`7�I��hɦ��J t�i��&$��*�$xB���ޓ�����7�E�X�4�W�֡4X��hK�I\�c�Ǉ��O���eң�cg[�E��pb;�e�uU�cA]pm�0-2�(���!�G����`<�Y�EA�,H���x���-��Z�0�Ƃe�臎��Z:��I����+W�����q�	D�K)����QT�i��AN>�P�����}j�!m�^�.)M���S;�^1�R���Y.��:&n�mږ�~�K�c���K">_u��nh��û�����tz�eFu��BlRH�����)��c�sG�X@F��`.;���7P��!����G����x?d�]���5>��Y�ܥ�FY8m��h��j	i&/W���4��aO]G%�a�k��a�D�M볡��$ޑ���(��J9��k����'�}�HS��9��=�x^���}���� f'��V�}�ނ ��΄X��2f��������tاw��E�k���y�k\_5ܹ3g뙘q����,%ئAW(
nܸ����je�N���{<���߇��~��n�[���W���GU�7��Vr��>����+<���97*/������Z��>����໻ܼ9�^�����������X������Nᴺ���e�q����!r(JE�3k=�?ړu��>\B��r�N0�R��ŀ"t��(2�,�oW����4�����s�If�р�7t]�wr� �3 �$7���J���gY�{>�e�>ж���'*�$��̒��K @����"��wa��!��iJ�t*It���'��E�u��������5�L���<���xTۥ�����
c�u]�הe�j��\�}��Q!���K��(У)}�cS�:�U\�^�$�??z�?��؂~��67x��K�j��S���}���M�}�ϰ�}���{T�Gmy�B%d�V�4A����n���S��W�w^9l۱9:�Z�p��5�i������3ކ�3ۭPm�-E��.�u��{|��,-�[#��g;+Zr��vE�"f8X�*vw��b��rCR��}�(����2��k�>E'i�Q��4}�O���T��{�&zj��$�"�a
}�"Ih�:�U$[{6X�q�ӣm��'b����Q�a���h�UB3�ApG��%S����@�Jj�4�i����8���M�� �����oJŭ!��q�<�{�a#�d�1),u#t�F�ګr꺥�"�YP�E�y�2g��|����O'ڪ�λ�3����5�7~:[�ch<�� ;V�ł�W�;G�=ك_���C�����ܟ��Z��Wa���'�wk�y!��_q�򎍉Ϋ�Oy�7�o�*�tk���-y��l����-�^�69�+_y�{�p�'�"�3��w�f�m�ͻS�Y��s}�>EQ���O��mے�q���bSc+��(�r�ӥ�[�:��^��������$�Y?v0��� �D
�@Щw|��NIr I��F����9&�?�J*z!q}���
�O3�p,k�� 4}P�wJB�;G�%*wX�F��"��>*��F��+�3��΂���8$�y)c��L�Kr������z�-���ǆ��X�!	���|ܗ3U>i�] I%r���)R�w��8-��@�8��f��z>'(�t�%]� ����]�.�u�y����(��V��Ag���l��(����$��A�@�4�aE���+T|A�B��]��υ;����c����x��N�W�%��d�1�X\�RB,�,v�޾�6��a��J���'|�Sϱ<�[[cF��9ܾݒd1[>::⩧</��";;{�Ư��ɽ�<��K���6�Z�z�T�a�Y��$���m�a�h��,<+ƃ��)%��+W��$!�B총L$!��CG�N�Yʬ���9��gT�}7\b�p�<4�e���g$��)�74�G���|\-�}�ŦONX�{��R��}dt��/x�UF��Np�`���"��+IVxF��ˡ��:E�j���H��p���z�s�t�����چ�}�k�X���܏���{��N$U�_��7o����X�����g��[k�+_�?����ί���Cx��i���4-W�0T��s�iʕ+��~�\;<`6���w�os|_��� �7��_�7ଙ��ks&	\Ia��񂮃jM���Bx9`L�y���샹y36q^��<��\���v�C�,/!!�˪X��wZk��Ğ�e����B�	��gP"]n��#v�M�(��P�쵮k&�f<��&3��]��Z��y���K�*�b�� !c�ܚ�,���\gc�
�����b�����"��z63�dj���P]�hc�"Σ<�8<�%�	M�0�;�4��\�W`�D&�u��:�������|M�b%��iܣb�u�dCʡg���c[���]6� �)�,����k{���)n��ܼ�d8i�h�!�����/z\�����9����	GgG�����j�$��vG��l�'�S�����vr~���_y�ɒ�Wn�9��p�+З?drs�K_���%ǧgk�zh}$p�|���̶�r������%*��IB�5�|̢�nK�Rl)F�p�H
\� ]k��0%�� 
{�<�o��t�k\�"T,Q�L|���M�&��QyT������7H[+@�~{��Έx�P1�)�ЙŘh�lTH�u���} �K�5�_�܁�	�Sl��&kʢ��س�3�U���b3�0�h���!6�q� �w(���7n�s�n��Nެ�����Z�!��|���;��^���ܴ�
	�sc
��s�կ��t�=�����S����o�[���������g�9�E�$shrh��M�C��7a�Aƿ4�&�&0>���?����ol)\}Y���2�����/*�j�'q�]�������$�;�������@h�J4�XVI$�S,Z���$��	V�f )1��,�����%�{I�X��RQ��:�>E���k[`=w��J�� �CP�18�e�Iu�"8�M�^�H=.ڞ-�y6����3;,X&n`c������ͦ)hip}��R"�B�� d�|&��8�V�#.%�*�͔B��Ћ�c���H�Q��48;�$��"f8��c7T�b<a~��[
fy����%&l�ͼ��8\�$�G���'H�Fȶ`$
�,�ޡe���+K�zrO�PW�*��B������(\S**YB@��iXU��/��꺣i�Ir��	]��"�|���캎�j�Ç9���_x�Ltt����V��Kt8�2)�JqrrB���7t�m��s�<��
cu�b{{�W^���{�8��E�UK��ݩ������rrr����׹{?6�Ľ "���a��?��ɯ,I���>3s��8�2�2�ƞ�����#�$�� BZ�� i'�?�?@;��тZ	�FZ��� �H��k5��~=TWUWUw8SD�`fZ|fv�Ͻ�}/����sN����}� _}����̹�w�ݬS���ucO����#_~�E��i8�͟�W<4��=g0����O�
�V�I��6\\4��8�:��&���Ȇ��nS�̡gG���>�D�ͶI��H.��3W��3��h�{�y�[��r�}�&n<4�=�Y����<o^�^5Gr��G��4�����/~�5� W��}�d'�����i�/��_�jK�����s����Kh�������(������Z������/���9������?��~���*�� ��]Q�w��|{�����������o����c���������F���xq��J������B�a��/�|��M䒐�8���홾^Uc�ݳa��^����7PӜ��Y�=����6�=M�Ę���!䌦>Du+
O&�R{^C�vVی��6��t�����?���B��Ƒ/.fM���Ӷp�SX��T�4b\���Ku$R|Z�P;��L��NYJ[������j;�G&�hZg�C/1n�.?�1:t��f���m%��������_���������f���1G٦���X{���m�w8|c��BKc��[��.؇go�p��g|�p����A��p����9�u�l�`�K�����{��o���n��~��^����G�⎿z;����gp}yƫx���@Ϸ�?!F����_|���cO�������O{�-��?;���q���-�~����zCG^~���?4|�6����k�����ဈ��7������?�������+��g4�8H`��O�xK���E�ύ秀X���/��{�V22�;=�^ps���'o�x���+h6p���{�)k㥏8���A�W]Ҏl$�<�>���%2y��aZC�q�L�����LHtt�b ;�8��Q���|0�a�ף��ȳ��ϻK���|��'�?�=����s��h/Fn=<������������7§/Uz���|��g���7��M�|���Z��������`~v�p����<߀�v؎q0\Z~��o\���5�����naz�����?�� ��;��|=���w�;����=66��oy���\��_q+��gA��6�#_���I�D?b���ѤfM�G%0k�������	YD-n���-��Y�A4�lc8x���0!j屠0H�7c�Jl�<T��%���D{�m��<�	��[��X������E�������x�ӔF��E�\X������iP����,���&b#O4��Fms>��6h�����D��"�5\5p����VUW��7�����4�X讠k4���+��?�s��{����o�ղ�`0҂��/������������5��.�A�ݧ M�0V�Q�$A���]����������_����s�����\<m�ru�g�o�utI�u�M��E=	�?ݚ��^ƤS6�|������������O�l4Hc�3Ʊ��N��?����6?�r�~��@���8$�C����A(������:~��_b�f��������|s�u��8���#l���=}�sq77*Y\1p<z�rYr�����=�����k����HHj��MF�I@4L���4F��m�qO9dRn-qw��1H�c���!�(�xFBP����M����!2�7b��5'=qR����ٰ�nٌG��������/�I�W[�o�Fǋ��O������ _=��<����g/�m�	۶Cx�����4��p�ϟ3x�*�G�G \�����7�|}�a����?�7�|ŕ��w�~�S��A9}�����ϓ�Ws��x�����8�����|�~�%�i��?9������'��?�35��@�[��w����?�cxq	_~��r�e�R�g��4��s�78y{��').�r�L��MT���M�g9N�\˖9�,����8�o��*<eU�|��D���ӟ��ׯ_s8�?�SF�����e&�2������K�m�@�1�v�-�BL�F�����F����Mo#Ah�bS񚠵?|�ж���K��h��^v�F����fg�4�q<��޴s�!�T�A^S��u8���~�����{��y��Y,L���61OV�T����}0�~���n<�a��-��9F�wǗ��w��=6�����g���y��[�Z�Hh	S�y4��37`�7���3Z�Q?񃛿��������g?��h���{z0�����_U���>{���Oi�@v ���������A�+�f��;ᓗ��~�|9x�̓�N���?���?�k8�8������������`C��&����#��oyu���a��zW�ㄓ@g����1I�������V�:��m*[׿��`_�?*�l�]�Y��m�N? ^�>E�0f�z���v�i`c,�մ�Mu_=c��F�o����3������&����Tx��E��p����x�Q6�0`�����;l��~�����E&Zz�̫�?��Ň����}F����p����E�U�W��=&\;~�ip?����������#��?a�lC�;�}�K�ܾ��G.�?AZ��~����{���y>a���8�5�^W��z��/����Q�4���^���[����������g���MԚ��s�I}#n����s!����^�8?��6�$k��:�W��!z��09B߰e�nUi�0`�Ehc�٨z����Wc���cJ�oe ��Aa�0q�0�����ٟ��/��)۪۪tʐ�V�}E���=}��nB������yǋ���Ep�L�tVU�.
4G.7l�(�?��R�v����<���/����W4펩SB��ۿ�lږ�E��	���|s{�����Ý���+��Kxh��~�M�]Gs�������ׯ���?�ѻv�Z"�a�\�n��g�^�>���6`��Av��A�w�s���H�$��{����+���3�Q#W�?gzx��A�i��WL~B�����9�/o�����-�n�����kB��Z���Q�-�O?��{�:���@?x������o�4xE���'�����_|�fs�_��f�tL�5��g��o|��N���>L���M<�y��5�������իW|��"f�w{l�r����m���-_��p����]��7�p��7ʭ�~����i��Cx�����FO�2�a�i��E��HG:�ʝFR�Նa�%�Ӑ<�8��8�G��:��C�rr��Ѷm�/�_�^T�W	M�mӾ�Y�fDtw�%G����k����?�2E#n��_��7ZW�MJ4m��]����g�&�{�ȱ�W ��\��z��p�vRQ'�����k.�����t�����Üy48����	ӝ`<D%�]�q}u�F��r��sܷ���>ph�i77�1�~��?��/^p8�ׇ���_�����v��>�2�m{	����6e5)�y�9����o�M-�&c۶�߿��a��q�$I3{���8'&�~��X�X��X���f,���iT��W�z�b�*VM��!�[��$��Z�dT�+�i��#�㈿�Q�����������gp��8�p�Ϊ�S۩�EH*��=�ڝJ�/_v�#�mSd`�$�����a�F���KrL��jh�����i�o_�
�0��W�3Bt4���x�qlyxH�s!������ߘ-Z~��/�+�i�J&~9y�_t�l���;��!�G��7X�w�4qb���f/4�?�\o���i��i��a�����5p!o���7o�۴|7\�[B�9�0hh��_�l6;�0���˿���O�K�������g~�󑡇�K����E-{���3�<\����;�y&�`c8=?z�-/�kFp��1C�3���v�D"S�"������a1o,�?0�[^$n�Z��?��[v��a
����[AdF5H�VW�6yc�N�dX*fN)�%���񀺚�0�gߦ������p����un6@�{�
oX��ӧ�n��op�=����O4]����������7�k	�"��x��a�v��m�B���\�,�WN�z$ɨ�W���Q�cTu��W)Ł�%o��U7�Q��0��9]Ru�)�n��-��n0������~⧿�c�W2͕����	����#����8�؏��űm.�V��Z��"�m�窖�"!焤ŧ@E=�6;�	@�7������ư�Z�N���C�ÜN z�!���x��=����hSR�Hr �Q�L �%���01D�D�FQ�$��F]hc���	#4���j��z��0�C �k
�㘐��8<���掮oi�m�f`�|{�zލ1B �gw-����=\���x��WuO�_��8�����~��^ r��~�o.	�/y5�哃G�����`�����?�nx����?���
�{����7q�s���R���v��8����:d���4=�7#��>�`E9�/H�1 �͆�	��������l^�?���ߍl6>�|���E#�޼y3�5�1���W?�&E�5#�����?��=Ӛ�c|�$Q��%_w�\�f��ie�ث��G/��=��\\�n0��+2N��s��|���H�=��6>y���|I�x��E~~L����H��T���[!�R�Rhyocr!k�"�S����hA�q[����e��ε6�/�}�E�r$�G..�ZdFa8�.�&�us<��\'u�$Y%O���p�������FU{0��8���w�p��Lۂ���܆g�JXM�?��K7�y�
��>�WuK�b����^��0���%���Ye�zL�ZMÜ�͘�y��������4�-S�S H�b�fbf��)��.��G�x<��SJv���F�{Hci�f�u�v$�'�ߟ<V��9�F��7�G����ZD%T��S��H�X�����ND[�r@D�'L#� �sY�8������������\]�Z�p���PUU�������k��-�Á���I9�D����1y�@�pw����W)B�^�{��w���?������������ �@�N���R��`<N`#�Q��nˮ{N�1�� ��l;qw�&n=?���{��q�ٲ���?L�����݅���0l�u� G��_�F$��c/�ƺ���]w��?m��:��q݈��x���}�ńT�̨���/´U��N6�3��}�%&�1�48눴�h�>�p�6R�a�'��iR�&`|�DA��		-�i�ӄͅN�&��!� �����Sb���C*�Ph!�0&�S������L��~r#�dՐ�*p���A�/��zEb�{�I8�~�>!#�ؖ�����1�w�1�;�G�x�h�c,�o�J6�t#��{!�&�"5�u�q�)���!��ސR7����A�rR�A7B KCkZ%�!
�(|}s�����?�[�-��Ϲ�~G�`��c���Zg	^�A���h���n����e�`�p:3	'N�e��{��h�7i�5�z����MjPXH��3�xћ�к9�M��@�Ğ�z�j&#^�A���	��Ҷ-�FոS<9}�Ec�)�ə&}w��sΝ�я��!6[�8���Ĕ>�ha"�;����T��7=�kxy��i��=A4�es����+h682�m���˖�����?�^4?dj��[F?�⧌�_e��+6�Gh���0��r~����<3�/'��0�qqq��+�G�^�Ks�)�+��n_���=�F����%��s���4��7�0�[^���i
�(�dz58Q�,�8�<�D�\�@מ��%e�s���<��o���l��{no5�p�	��`���1*��=1��r�rDS�<�.v��M�y7ͷsww`0�wF�)G�1��#u���|���*�g�/I�;/"�8����k"�9��n�]���(O�6��77G^�� �����%qv�)�����������x�� K�NȄHf���'E(θ�c��H*r�]aRi2R���A!%8�Lad����D3&)L�0��6���9c��mdܿRx4�J,��q=�5)J\%�W�n���B
�6����c�OZh�����m�� �r��$�&IA��10ۻB�>BR5�)\��&InS�te���ن�$��3N��O�ُ��;3��lP��$	�����B�g��� ��~Ř�Wo�M'l��ֶ�)��wF�{�#���}&у���轐��m�ѵo��O~�y�s��w��{R 1�6��&ڪ-�9|�D}��A��4\�Z�j����2C���+|� #�L��B���kp`�C?p��ܴ���7�����?}��^�������/�;6�/��oq�;~�S��#v��~��?<pu0�c�h���[Û0��#[�dnC�1�� L���5���Ll��e�4i
���l�j~�W�g��>~ˍ�i��2&���+��7]
.I�7!�A0�M0Ljpl}� �G�ǀ79�*�8_(M�eǌ���u9����˘��Ϭ�!���g��Z��r���wA.�u����14�i��1��){���8!�����w�H�t4�A�Q��!"2��wI=0�I*#��9�)�䋚h�ȩ�ttJ���u��Y��d��Y�~&��[�	��|1s�06�m�V=1��IL3Ept�p�k�|{O?�d��S�����؞�7�b3����\M6�e:O۟�.(.	��>�ǩ��n�6��#QĜ����j��zZ���SJcR�T��1�]���2�O:��4E�7�(&%sK.��!uw���߇�!1A!q�af@�wd���c�u�C�7��v b�ڧ�T�p3x��!./a�i��#����B��ݮe��o(���Ln$�_�������˯��1(n�>��%�0>D��H?�SeM�l�SC���p`.	��I�Y�K�#$������{�S�mk���M{=wwo�jU����3ǫW{��&�����c��rF�~b�d��2�{���z^���[�R6pq�az�>2ӥJz�	h���Q׮��H#7M�V�`��}8�K�">����'qWDp��E�~H��V��M��c�����>���Hy6��x砜�<~N����e���oOĥ*��B�?�f�L�:W5��|0Y�!0e��� s��T��:6ɶ����u\Ȫ"s�������x1䵸�"��=�<���c޻��1�T#uT�!K��<�FB<jFEg�x�r��k�����́/��m��KKg?W���Ѷ��$8��I�iF-�X�?D=Ǧif�*����@%��ҕ��d��6��|�
��&���	1"�*���'��]J�������3פf~?��h9&bT��a
?I""B}Z��a*�0��T���䬢��^~1���u�M��!��c#"���ژ�X���B n���[ڶI�,���&3Yj����-WWWz�f���W�~�c~�ŉ`5>I�UP��4(ɞ��)��ar!~���#o�>�~�ߴ�#��z`�q�fR����\]/�.�����.��~��a `�~�	Ǜ;��=bq�臟�=���4��p���]n0ہQ�Lt�i|�w���|��߀}o�`2�r���n|rU�x��ı4'�4�^���=>e���⠁ ��#&d�=Q�X�3����L"u�I�gg#ɀs �P�N,�"�vF
g�$&o��In�%q�!#����t"�0��H����rz�삛C�mZ#�t 6�Xl01�腽��)��U��9�5���\'�mҷ�HTk�HT�ֺ&��(��,���D�{�4�I��Ebb�������<cB�]kd����0ݣ��'5��ݎ�1�v{v���~�_��?�����\\)�Ȱ6k��lMBʅjN�y2�B�,e���ly:�G����"��p�.�w��d�qQ���]E�k&�mb>2�1Ib:��D���§���>!���$��9I
Y���9p-�ۤ��P��F��������:�pN�e��{�a߶F�4���n��5Z	M�ӵ�������d�ā�����w��@�~�7���ɏ���̐E&�	�7,�Nn��o�O�g�����$�QYg�������xdJ��-2��dN-+�b�����^�%ƘD5���T�uyy��w�����g3w{u�e��]www�ݍ|�e��Rl��5�u���o�����Gˏ����A.9����~r���'��0�|6q�`8:�7�	��ah��g���M�AR���7Dq8�����*"���76!�tq���F-����Tb�s47�����ʏ��t���m�s���_�)��宙�����'dM}:�mU��`��[B0��Z�$�{���p�4�M��tM�Sb�tH�%�M9)#Z���4�$	�g�9C�����^��F�mSZ�"}g�!\������5 ���i���i4��@�WuO�!�t7��ϟ3����z�={��0A=NĜ���+I�i�s˼�U}b�U�V��P��cV�i���g�������f��Y#��`@7{w��8���2����R:�M����DN:�Y*���RM��ϑ�C" ��s�.�o6��X't��x�˫+vێ��3.�q�M�I���iPo:И��:���O>������;Bz^ډ�s�&��|�0(Ñ�j�۲1W�C�o���n��g>��e���|��H�~�6Ѷ�G��&��K~��ۯ���ٞ�:�p��+��0���7|��xn<�QS�N��t��tx×��|����oo����K�է|{�-7w^~��׊ԼV�2o�`�;_x��x��=��vϷ��xs�ɲno,�d�A9"��g`M���o5C�.�-�m�x�b�;��/�ާ�á���&�_F50[+����&�T��W:[�c��D�������āG�]�J�.��:x?Ɛ�c?�7��<�1��+�������8�YR2��Y�gL�H��=��H����:>���+�v{�@�Z�< �Xi�ƞ�x�s�ttN�p��i$d��6M��C�,�Ѷ�L܌�M�:�1�D"���D՗��l6���5�_�r���~���B��o���|�f�����+w�?���C����+��C#����l��sw��04�ƀ��m��{e��G�;p�I��4�X�4ᇉ~���rV%���=�6�=!Ll�Wl��״VT���zaLI�H�����c��p��g��N�p�s!�b1�{2<�0q8�sk����Ξ�Y�d���)�#@��4�ı7>}�Ǚ#�ׄ�qL�7ӑ�5�O�;��4���kO�z�b��^�k�zCr����͝�^����W/;����&��|y�~�՟����	��o���<�X�8�����3�=6���Y�|xx��'*㙑��ȶ�-�������w�w���+�����o߾�a�mf�n�Q��#����$��on��W7�tQD�,E~'�俢�Y|g_�h	�cLG㶌�9Yv��͏d}c��v�x��óg[�?�0>��p�v��m��fU1x��G|ڳT�^?v�Z���~8�U>����X�u��n[�(�s��Sr��!�tCr�̞9�K	!�k�����k�o~/�z�٦\��%���v���l:��Zw!�B}�8��q<S|F�r�\����/a2q�i�t��8��%ad3�g>�i�,A�8�.�#&�C��u�����"����v��|��%"���ӱ'G��
ZӠ���ܦ�[�v^�*��:�u#����J�p=���h V��I�gn"˞h*фq�ډc��t���N6�m����x�H��n�I��)�@D��I�-b������f]�\�-F��xd�z�ab���~�4�|~6��6��K��iL����E��:��#>ݷI�DV�:'����uן\�}��G�	��p��&b���%k8�Hs%|��?��� ���	a����u�}�?��Vq���/_ꝋ����_~0v��#}oZ��SC��:�:�F���;����O�a�&���L	#�n�l^c����cƻ?������ô-_|ḿ}�'��ᛯ5���6��ӆ�lE�#��"��t�=��3h>e�������!p<D��"�V��ӗ��������}��F�x����>��'*���S5��w��b��~'uK������o��04-\m�T��p���}�p�s��S��O�{��X�h������!&���8}��Q�1���\VӀ`�H��ɬ.�}{<���O(!;w�$[�tR!�j�B ��f�8l#϶\�0<<|��5����s��?�&p{{��7tQ][�pu���[����1��[��a:�x?*C��OD+Iqc�0�vF(�Hef��~����������aM���5q�����ډM"��3����y�=!D�+���'cg�HE87!��6����0��qtL�7�#���^�Kc��}ޫ+���>��sRey�q�F�q��&���=�Z&k��)k->�Fr�����M�b�Çc�V��?螥��&1�O����V�d��k��?�Q������-֧`�	k�4����$��J�1���靁�nb�,S�9�G�� h6�Q�q�Ic`�d��c��Po�"�(��p��?���HR.!l��������?�}������~�=ގ3��1>H��H��k�#��?�?Ŭ����g�}����z�
�=�d��ܹA�57�+���\���؄�������kڶ���ҵ9~�ЏD�s���������^\cv�|�qox������ݛ#�7=��<����3��.��}����a���!Ju��H��{���r�$�0�Ol�!��i���t�a��3�����;�{c$�J�&@+�Ĥ�N���b͘9����X3�	2�]tc�i����wȕ�B�Қ���8^{�ه�w�1�17K19H+��"@c�UU����O���v��i�����Ȯ��vj�Ǒn�b���WێϿ���_}��~�?�eF�jka�;�>y�h�ؾ���dymM�h��5Mt�����݆!$�q�Ҷm�{��9jʽ���R-֤v�Pbbb@ئ���삪��5�\��N�jw�]�;�<�do.�1���HK�9-EVoi�r���W�z�W@F@�q��Vbd=]'��S���J�u��s�[1*"wN�n��n(��9xR��F���&�����0�l��ˎ���0���Q�̶���+�&�d���})�JVSOL5p���{�� �����7�7�ۿ�`���Px�}����>�´��[�t�8��w"�&�?&����rH��!hL��������p|uGl7���L���'t�;n��0��:,n�b<�#q��v"�[���W��g�����p/�4���%�����`w��v䡿K��E]ʢ�R�)��Q�|��`��>0ى���(��!�}�*�L��s�5�e2z�& ��D��m�u��zy"{A����f�Y���"0e�ǘ}���8s�R
f�V���y�%�UH1�mV�1�(�L��N��!�q�y�>��O�1͖i�qb:<`vk�dy���r�혎��/麎W�<�ݎ�WE���t�?q�7 ����bMCR��6;E���Ș%&#c��Dt��vO?���D�U��AC��|s�����8C��[\�#�Ѯ��1�C�.�x|�@Z@a�Z�I�F����=WrA�6�d�F 7�S#��
>s�� ����oq�Mv�N2�//m�OQ١po5�?T�Eʃ?�>%0Y{h9�.���6L�h�L��a
=1�^h2���D4h<�0��g[Lr��I9��Q5N��qI��OI�|Q<$Q�i�W6BJA"��DT�1�:�I�1��aGC���#�A�=����Ö����i������ϳ�����0��
K�̵����v��Ա��鮯�M���k��0��f���X�)��a�p�͚���sp�G^��#����,-��g������Zc1Φ9ir�a�3w������+v�#�����'��Ef��5W}k�c B��dh\���:�IQ�G��p`�M�Jbf�H�����{�}3%ik�:����I��:�����?��!%�j?E�Q�m�m��x9q{������!��I�1yO���u�k�D���[�_>$�#��Ֆ�E���#[Fk��D9닋...4E@�suu���㐼~L��'���
��&U1���e�k�l#&G�&��Ügj���i���ܼ1q6���b�ڶ����&WQ���dK�k�p�4�6U���~�8�`��ç ����n4} ��%#��N6b��Z?۪�ԧ6?K=�����"��%��&�V �.�˜o��!�IYXsne����˫�)����C�o�$�x�aW#��w٨L��N�-�:gf����~�����9"��4"�#1B���J�iR����ߜ0��t�,�����'�w�ofO���oy�t8`;˱̹��GA�q���}����%W�7��VF��K��[x���ޘf��czp{Dn�õ�m���0n9������5�����[�N���:��l�A�?�l�E%۽�1q��ǔ"��hq���>0{-�"v$�7)����^ъ��s5���z�g<����]�Ҵ[6nĴ�+p�1��1ıg��Ӹ@#(b�v�F��Њņc� ��
����5!�(��*CKq���� ��T�@��c�j �9�R� ���ѽ��,]�sW�8�븖*�l�3I�5�z4]^:nn�v�����5!z\v�k-��J<���ֲi>
�� �vH6d�ߤz����IW�bƩ�͈�a=�LQ�њ�R;.p�1����4mæ��p�FA�`D���~��`F-�g�2M���Ar����� �	Ќ.:J����Y-�3�9��-�s/%���x��0�'�
T���u�{�X��&�ߤPu\��D �Xl�8�I�����?�sc���CBvδ�X	7��`�83.�t���LfF��@0���:�Q�9zHj�d50>���a���t��.�2"D1p��s���¥�LX&�D�t#��`G�e϶`>��m9<l��o̋O��[o^�|�e?�T��}����7���/^�������g��)"��0������A+Nu�C��5�7zX�~�i�d_Ѵ�06��G�V��{��;M��G�����)BRu�W��L��Ʋ�\3�-�WWW����)�(�1�6�9H�b�m��0L�ɗ����I~�ֶ��"f��?m�/,�H�҃&j��	�1d�s�@��K���GMnABR��Z��'=|�!���z� $d��g�w�n�i�᠞������l6��s�����@�q�^��9�[��ǁq�l���p+��иbD��'8&��%�ўE�;6�U���ȔJ�Y����jp�0�Z��-�Gг�a�%ަi��Tc��OM�a��c;�m�ul7]��$�w�y�G�����Y�h�&%�l6�6�9�����6����x�cJ?p��T*Kc� @����1FƄ�7�M����إ6z^.����i�hR�19�7���M�8gG����Z�Z�$	$���ԫi�S�J��4��s�8�j�B���s�'��Tߣ��M�A�M[�&*QQ�mw�Q�yE��L\躓g�����k4�����9�L%�NN	
?T�(H��1��������|���[��s����ߢ��?���ȥm���pGG��15B����q��o�"0���Y�w���$�8xO�t|3�+�l� b�J�����f�}��p&�q�JXa`3�A�@H��>L���5و��O!&�y��{'B��1���v�!��_b��?F��FdH�t`� ���l��&W�ƣ�a`�'��txP�b��a��#!<�kn[�@� �l��⣦"h����=�-4a��rv������BLa���S�#G}�8Q�T�!� xD"�����g_���>bLO��8iE��F��ҷ	���c��ن��р�˫�X�1�4j����FE�iԴ�ưi�:�i"���l�{|�� vC�g�cS3"���x�8h.F"=���H�n�lq� )2�v�-�6D�"[������zp�\"_�80\�����6'b;ϯ��#�Aj�S�*�\
s�����o
�&UٔQ�>Dz��"��-��j��E#��'FXܺ��<0�*4CL���A���V�ڍa
��$D-"��ӥ�:xy�fG�I�L^;C�.��ع-�����v�8���0��v��n�	i_ ���{����QCi��@wG0W&�������3��7��:a#�FF?ll��A�ϟ?���O~�v�����ϟ�#����ꊭDd�54u�jz��%/vo9�X��vt]Ǯ���ϱ�h�RD��GQ�oQ���s���t� \�=>�#L������H?F�4���O�@�"���s�+�O鐁Ș(x
��H?�D����빳���{����o{��A���a|L�4K��G"-&z�#8!��H9S(`�MR��^@!qD�{�!�i�TBY�Ϯ�bJN��)$7�锂��+��'��r��|,i�"��i47����L��v�wb���#�L��(.���q�����Ns��26���k�ip�DKO�qQS[�4��,8��,�E3K
�wS����v�*��6BHU�d���5�u�vO6���ilU�Lg��}8��8�Y-T�2�Bvw�k�%�$�2��ؙX�]��R�ue>�G�9��d�#�I�sy��������#2�&�J�76�!�����4W��IUf�Ꝛ�X�)v�yտ��CH�E���e�x���f�1�(��� �n�E������w���P`z|�c�As�Z�?��C�?x��?\���C0#��X�l��*	x3i�f�A��.�v?B.~�C��i���QD}����	`2R��nʏN�UC�R��CO�<7I�#�C%�ϹPb�c��xv���1�<�3��(��:��('d��M1WQB׏L~HȲ'����Gr
�=��\�&>@x��{��83b�#�O�����x &=s����:�$N�@�ؤ�D:5��G&�a�_2���(�0�r�9�Lq��>x�Ɵ�H�����	a¸��WOJfR�dC��,+��$ӄ�BkZ�O��[�xI�M8��b'��#�{��k������F?��Z����H��� F̜�9��*�#>�3��1�G�\�7��C?#�e���YAl3�U8�,�)�Q��D�K��cN�p��g�A��.K�e$ŨhZ�#��ϕ ��4MR�y�q����H����	k,mץya�R��HcG����c�P6^�&U�G���n��ߪ���TWN�) �Iu���&�h��W�VFČ�>I�. mqO�{/~�6�{p{����	l������Y�h��8��q�e�fh:G�&�{�h�b]K4#b��<�p�Q��խk�CL�����sʟ��0�i"�0s8Z�'qI��En��eS&�g�c���E�8�"`MR	xB�@מG.!���D$U�������'%A#����4$��%s�#q��~����A�q��#a����0�bS.	�o	j����7��3'��~����5f?u�?�8�WcY(\�������"�e�nx�	�#��3�'��a�99� �{e����}���<�9ce:�è�e�<�00�c*���]'�u�3kd's�H��aiVm�S&��[���l�̿w9b6ݹ����,�ٞ�㘲���\����/[�ˌ\�{�mW�{K�%�ID��;� NR�IZ�{T���#!ݟ2�hy޳')^(�j����F��k�V�26�U��zkIg�g%#���0�4�.�UIpa�I�궝�4'�8�_Cn �'����4Mq��#�.�tAz�ݱG���Z�A�%�I]?n��k��;�q@5����U��
�II�cܩ�or4a��/��N��	���K��3 Ɯz %ފ��r��L��9�Ĉ�  	�!Q��rQ��euA�dI�~�X�i2��Y�P�^`2����e�1]��F0]R�x�.]���2] �\eD�c�S�t8 a�O=��`�5<}���#��#�[\w�5��k��b����~ĉ��.:5�bwD��`�`a�
v�?`���qw�0�d�t��rF��1�)!���m��&'@;�Ê��+���s��xN�s�H�Bᔲ��>@m"�D�����'��S] ��i�#��O�BC��}�����/[Vk��3����{O�F�h�?I�Q�G��l��A�} #�ܝ��{T0%�;gJ��3�c�x^�]%��ݕS:��L��3B\�hl���9�0�f7�ƇG����5��5� ��(<��֎-}�)`��������1�7�hp�ER���$��Y���Z,��l	��."�@���&|8b��4���/qW��Ն�!b����)S�z�� jE���9�	�.^�Լ+C��fv�Y���9�9Q[�s4e���r�]���C�w򨩬%��� ��س%�]�Y���o�k&���#���d�g�Mp� 3�S���w�矾�/���!�ݷ��
8D�� N������Q�#1�3�Ǐ\��bD觃r��#޷X�!x|T?��:�i��q4b���3l�MJ��a�+�	D�g�/���I���	%�jJ0皜g?�9���,�v㹤�s������uѨk�5 �R����Q�z.<��>s�wEܭ��ϭ�C�Ϸ�DV����1z�}���2���*aA9h�x]8��fd�%�s�9�ܬ��Qڦ8#R����=��.�P�W�K]nS�����9»�-�c6�S�9�����f�	B���:�g1H(�	ɕ�ܬ1(%���YLw<�1��C��ƥ٩7��:����g]�����߷}�M:ī�Κg'�Si1���h�Գ4u���H�GC�:dj!z|���H2����J�WKg��]/G���=>����8��<st1��j�N��$F<��.6��'�E=AT��Ĩ@1���9�T$�e�Q���i E��!B7�?����$�I�Ӝ�%�����*�Z�4��9���H9�ldn��!��X���M*;���8��@#�)<��#�[wL�+�p�~��-�;�Sx�hF��1���-�"h/��Z���Kc  SC;^AT06��5YsZ����m�C��K��;ߓ���ESܹ*%��Pަs��bE�d� �
�\7��F��3IMN �U4%-mBƞ`�1�̈-�5��򳙠��n���(��SH?ƈMH�ܻ關���)pvP(�B&t�j�fn��Ǚ��d������ُ��+��'��[l����8���	V"�v�Q��o:FRN�jL�=5�7t���
������~
n��&�p��$��h��`�o��^#���o��!�GA����3������o�I�:J�V}�����-wBdR��'q��T�{��WM��ٷ5��ZȾ�'*�[�H�{!�9{����r`%�svĜs@����O���ٸ�x����Yz{d�쒓,/n�`�91�oZ��u�h���V���Mk�j���F����1[��e����iSó�+Fo�L���f/?��R���8y�1 U�͙+'�j�\p�)9�y~^�υU�3ɲFz!�$5��i�p�/c4|_�?���������r��3�*�R�aaH�`˾�s_S�f��St���~rn�y����x}.��D�gg0&2{Re��R���I	,��(�5�ë��hs�Ҟ���9���v��6XB�{޶-��0L�!9�QRM%�NER9�m�lh�m��]�G]�m/ |F7D^�x��k������>�<A�J�8���rp�D�#�b�M�="v NGL�|��Uwj"qX1�Ns�<�5o��J���F��@h9`̀�6����@C��S�9�9�0��tRŤ��$�R��AD��1�{�B��S���l�G��͉��w�;��s�ٌ�N��|�(�������͗*#o��/��u)�D�x?��0z͕��w�s�G�n�>x�1L�C�,�k�<��:G����{I�@&����`�A���1�\�Q��F�pI�1L��dvZ!kG��0J �@�0�D"Zu;`�A�hDsLI����q��m ��(y�pV��Fc	~�hU�B$�l�3����9&�ψ2�HL6��I�c�b�9C�96b�Q �DR�DJ&�K$�M�j�Q�0�
���?��=M��gD�\4��~
j�,�Ĭ�Is�Y]�S9���S��	�Oܽ�F�8bc$������!�)M���:*�q�
�@#�Ld�8�S���~;qh�.x�m�;d#���l���N�kC������^�mK���䖛�DM7���m�Z�44�,Ǽ�i��a�����6=^��.>0����;����]�S~bL�������1Q9�����msΎǠ�y�Z�ed��質�k*�]�;������K�����.�sK9=P9�L��ye�������zt�ϟ��~v�7�y�х�yC��ӻ����qF��Y����-�3?�낄��Q�1��c/��ѫ�Z�<��܎�������ɕ��$����[�_ã<:�sx+�Y�o�g)M���o~�������3%a(��&��0'6����xi8�/R_�i���#��<ߜ��\�)&5��d��c��;8��؇h�[�q2bݨn{�&��H���5�2��� ���h�e�DU�X��o�v�#2I��ɥ��ņZ���Q�=��@7����AkB�?�K:���P�@� �B ��%�Ji�J�8;I��X$,˗M�|g��y��<`h��O��d�r%E���ɛE���&]A���C
�7�I�(�[��x�,!e/�Q�9�k4g�ob��oz~����� ��iCDX3�ޏ�RQJRd@��d�HرSwVc�F��~�<KN�+��g&A/1�y:�V�"D�D$��h����^q��8��@��4I�K:�9�}J��MR��`1X$&/=���$�`TY1��	>D"&.�1�3�%�ʞc&y��#��;!�Z%��-Ցpnp�AΞ��=����EA@\zR��)C��vϬ�^9y�s	(3Z9Q�L'��	�x��Ȏ�18�! ���k���Iwcݜ��a����8b5}���+���,n�����ih�\�q�}ㄗ�b7#v���D~�ox>��J�!��9���>���c�� ��t����[k�ٍ.]����2���s.��y<��Z;�Q��b�ϥ>ָ۳yU\N�N��.�WBs���/Y8�ٚ�ﳑ�}1�׿�}��Q�'�����B@R(֗aI�,I 3y�f��|��=_��J�$��Z��g��{=��������!���5.����w��԰�%�xRj-$��9�I+��OP�^���O��;j
���l<�� E�J*K��dM�y1���s�S�+�w�{�0�^�)�t~�_��������#"}4�����"��jp����&h�I,�� Tg-���ZYI�x���<�0SzE�:����gb̅�5�dh�ς[J�B�+.�9]�l��&�
���V�'�S�	/f�����	:�$r6.pJ�e6����/���NĹ�Js67/N9�R��h��D�x5�{**ድcp�p���E"��F*�'do��N�yH�t�h��QI�j}ڈQi����B�d��{��[�JBN���Ҿ�=G.n:q�&���ܟ3dcP=t���p1�� �I�XB�oz�|vM��4���AwgiQP6)Sj�T��c���fR{M��ͬ~PxV��천�W�B"�"'�#�t�'����9׌�-��YyZc��BTuM�Y��@��Jz)VM� (ވA��1G�i�C06�83b�t�ٞ�k.
&^a�e�[�0���#j�ӂ�Dbn�ރ���u��D�#&��m��@|��Q9�Sf=�^�1����0h*������om����c}��i��c�<�X�H�g�8���rJ�ڳKRFͽ�k�%.�� �������إI�_�"WP)Z��N�q�@�aa�j3�{X��P#d�>Kn%�.�0kD�?O���<���$�s��ZS\&y.5R\�&���8�r.���8_W��w]���W�w�ޫ�*uҵcTF�Z[>�z�������y����������01�#��.;B
XsF�x���H-}U���1'��!���h/�}�GC��eOp��	9��x�X�0#e��osC���2�R�r�'
L�A��A4R���<ŉ Q&�hޗԒ?����
9!E�f�DH��t�6q����L2ՙK���	��2�JTO,A���%���D���Z߼�DCH.�:��x2l�r>�=%�.FSG�$���ECL�X	4>{���$�	�?����\�Q�S���ٗ�����r��O���-�;��9O�}�Dx@���k����7W�̹y�9�1�v��)9��Z9ؔ�F��,���N#��݈�� ���Ѡ=㬊<�I$��Kp��M�*�ߒ8m��)�B�)�������t]8sխ�$ی	LNd�:������sҹLTD�����O�,����"�ؓ�!F���N?I���Rѐ%F]�
Vȩ�%�^��4�w|� �a�[�m�̎0����9�;Z�	�	2@��S|@Dh�%>zl�D;"��` B�`D��J�0H�6��!baj0��5���/X��Q���������r҇�R��!��#��9�4�N�6%�	Ʌ1sP��k-&��Z�6_�3��i��1��X���],=W��kC��_ϩ�4˶&��&C�����{)[R�H1?S�ʱϼM��#��*�U�L|ָH���R�]d�x�Y�\�G=�o��]��r_ٸ[�]���9�$�s�sI:X�n�gk	�Z��1�<��Kr=���-��i����$��ZB�[�Ίyt��{s��l?��N�]g���xK3�;y�e�<5���a-9���E�Yl=��xvw>d�hH?Nf����t�ǁq���3�����0���m�2�����r��1v�`��Q�1#M�b�W���y�i��b;3�����@��F���6�n1rvy���,�E`"r2��s��+$NE��6y�d�\��|H��������y����!Qo�HL'� J�ѣܒI^>�ԹF�_6�N]+Wy���2���bg�,�1�K��X�����SĤ��N��Wz����#FbhQ�|R���0Z��=1h@X0Zl�t6��b$N!F�V�V�~Ě�_2җ�y����f�R�ڕ�y��U�L)�夙!d���x<CB9�� �r�+�bɌS�g�s���X�z5X&I{�,�0�J�H��s�z9�
���� �F?"i%��s({��<��K�Gh��S��JW������[9x�6n>k`����$�	^�u�,^`������˛��F���#�`sAsh1�%�~��q�GD^ �1D��h�1�'��	��A�<�5�[�E�h&�M�_a�=�	�����S>l���^EˀU�rg �[�{I�k���S_;�%^kK^K���޷��і�m���K[�@��Y��Z�ε5���u.����8���R�=S���8�%4�,�+��5���~�����c�斿������9����T9�rM����O���3��Y�Y?�$��J=~�����L��{k�{j���eo�������k+��8K�x���Q�w��y.]�����ჲ��O��5Z��f�%9-�>��-C���� Z�j>�d��@��g��[��O�А�=v�j�9�#�w!��� �F`Έd�|�G��ЮͥF�KϽk�־��ez���rOͻk���s���"r��R���軴�z�KH����+Ϸ��vk.	�r[��Fl�jK��>�C�\��%���-��v�����܇l��ӏ#2!zZ�45(`0Ҟ�l�H�M$���`�A��Aӈ�5`[��H�9B������$����Z;�2>T����9������	�TUDʇSP�ʽ�j�?&rFQ�� ޅH�.���
�?Ֆ��<�������X{f�������f���[}nks�9�w	��k[J�T,�D�W�u�c\z~��-|~wi��8�,-�Y�Q���^�c.��{�Խ*�w���T[��%�3�aDLN�q~�6%f���BH*:���J�q�g�����0�6���#{�4�c�����f���vW��s}NA�a����`�LZ�5��cqd59��DN�*�y�i	'jM�0
=x�kD�lk�D6k�l�""�8K�bI*X������ƥ���"���R4������>�!�r~�����./��4�F�ڻ���_B8K�/��w��_C�kk�϶\�����L亴\ѧ`i��1C�8�f)�i|HD�,�[�p��ef&Sr府	8�AqJs L!�q���Z�l�rC�o�X-�C�ċ����KO�4�	��DkJF漓�S8���/s]�@"������pd�'��ր|�",]��Eu�K��Z��-����`�Z�ڳ%��S{�4�_彥u�ȫ|��)T����2�f��Y�UI�ʹ.I.�����F��Ky�˹��������\��JK��kgU?W����>[c>��G���U��=��['H�ę���)2���P�+�����^��|��ѐ�V �0F��R-c��`s���]�37рu�X�X�-�Q�0&%T+��I�N��1GF��1�/D��e����)��W�R�~���8���%@�9�����q�pn�>�i��u��՜dm�|jOqskb�n�䟏\h��<�"D���&LKȲ�G���$PYe�'K���]����T?u_K��c���R�?�Ь�y��a���?˹��kZK4L!�@�s`�[���S}K�~\�h���A3-5��v�� 8ͨ�5>�-DSS=���
}����yN�3��]1���L�Dfq'�-�=�W��b�q������ ���Җ�<J����)���c	Հ�4ǵ��q��<g��x�뼄Xj���bw=��z�>���Uu�u,�R��z��ޕ?����_�ʈॾkDY�p�?K}����?���� ��|�u�u�f��>�u��>�w�<��s)�+��ѻxA�	D�;��M.�Z�Q�r�aM���Z�K�IJ/�B�����W�8̯	ҷ��2�Q�Ӌ?�b Ĝ��%��b�6؆qh�b�*�÷s�5���e4Xb�":�p~A��gՉJ��}�~��zg]��f�{�w͙>e�x
1���Y�GN�[�[ز�k�9�%�FY
/G����q|�rY�C���� #��y�?[B�M�<����1�}���0����ٗ{\�Y���~W䔠0�8�,!��].vR�A=��_�~i%��-�e�6M��{&�?βkd��eU����Ѯ�*�"?7�#�͆i���S.5�6��a�8��tD�)����~��Gۥ2��J�{| x�E�����H@$e����?"b1�c�Q+����{'\L�[j�2��A��/��Ü��_unh	D��;�l�5�sz���Z��ͭ�jN�F���%���<��a(�Y�Tk���p�Kc�c���}��1�Q��97#��S~��Zϥ$X%1(�\kK��f&��l�`p	�խ���@�R�I&�OE�>%�,��&5��ǌ�Z$�IPs[B��3���ߛ��x<�k��=M4��L&��Vv��g��4�4!��ն`����N�}��ZnZ���x�_�}T���I%As���������*����z�Ÿ��(���ӥɅ׏���ǘ�ޜk����s]Bv�;����.x�Y�^}9�8�z�������\곞o�`��3�׵4�����2>u�K$����W�Is����j܌�K�&�Y�X�%$V�qi��y�{��s�r�]{/�D���,y�-�'�Ws��{�Z�|[���F�lΝ��=�w��W]�$E�F<�q��RbHp���8�m�;��b���^��Il���	&���0��#b��I#R6X��E��΋g�wm�{'�5�l�� �)K��0̔5��9�2�J&@�/.��S�Ļ�_BPe+���!���Xs
�R.��滄�r�E��K�ǯ�T{�d��Z�^s�K�	�:��y�1��������Ҝ2�YZo���:�R��V#�58�[=�zܥ�KD����>ci�K��5��I��._�D�^s	7�9�m��Y1�Jεd$i��+�aM�Øj ���	����{y^�9��i�?`���Y�8;xr�yAOp4�);U�}�a	b�Q�Xk�h������f�1�V#G�����|���"R��O�w���˽��]��lO�c��ғ��u4��~�H��K�8�汴�g��K�}ާ���,�E2jV�YF����(٧���h��n��/ֻ���mK�4���-�k�w��oq��/��)B�R��y²��"1�b��!�a$FO�Fe	��8���; @4t�K�	�0��_'�s�Ɏh7��`����g�&ep�u),*��	��B�J����S��w
S6�pD"3�_~^l�,��ZK��d��J{nq�5�!�Vs���z�ŗW�멋����r���H9�<�r���D�����j�Rr�O�=��N�4��^g���)5,!��_=�5��y,�%��Ԗ�����X�z-O��F��=���g^���x\��֟
�+�X�Sa;C��b4��8{u�ӄ%��U�?I9|�#U-���8�O����C�����J�$��A�yg%�Gb|:���5-^ _�B�*"��V@k��$!���4q"1>��K�t�Ϧ��)TȦnK(?_"��X�!��"�Hi�z���w�X��F�K�-�7?�w�*���tfK\~��N\a��q�
�R�@�o)�|v���(�}|j��E���jX+�X#�Kk^B��{5s���f���;�4ǵ�S��#8��}T����ŀ����8�Hd�q쉱�m��ZF�%k��&�82&"�=>�MR�R��jT���dh"�S27�3��A�G˲��μ�� J�?�t�%^⢖.i�����=/|��~���KYS�՜q�M.qZ5�Z��%)`q�y���g�%�\N^[g�K\ڟ�,��إ5�j�z=eĲocL�|欯�[������F����`c�yX�՚�+9�r������u�{�ϔ�y~e��᥆��߻�kI�X[��X�ԕ�^��6K(�*���9�� %����~�Ԯ�mS��,����3M'8�K1����P�q�����ؘ	��8NHl!�Ą�8bp��;DL�	LDF�DL�1N/	�M�5�����қ#!�iD|�ňФ���vx�1����D���p~��2p�Z!L'�o��X�<�1��b)�^�%�CDP�b��V�d�$��؄���X^��-���_��;���%����R�0�)	��Ϊ�=dѼ�C�hJ��<�z5b)�Ľ�{Q�����F��~����^"������m�1JbB��TI�ʽ�`�޿2Y^M��}	!媗�QK@�ϴ&����㣵����Ӷ홣FyN1Ƴ���j�#�}0�<&�.c��0�Ac}�@���8q��战�0��^�FcF�t`��4?q"LG�1��+D�c$��������_��ưϏ���C��Zt�1ƹ@DL�K Yi��$�q����,3#y�����Y9n��]�wQ�q��xj���kb��c�A�jUJMԌq�w���x����)�s_#���5׻���c�E5�S���k{�F��ߵ��2sP�����<���k���F�eE��K{Z�w��{�י�z���������˥������x��K0�_f���~v���N1�ˁ����b<�E���cI��>�}56�Kv�����0�<sA1j��P'��:���hiq,1ڤ���rZ[���ڶZJ$�jF�f�6`D�����:�w#������Z��|���ֈ�r]�8�g5B[C��K�ui��ƞ�Y�$bK믥�z��y�}�k[C|����y��|g�5�ϕ�+K���O1!�3�ڣF��w�S}%a��d��/���.�/�ԧ�S��Y�r�!��	~:�ʦ��ݘ�@����8W�3�`��:����c<)��u:���I��MS��H�&��GE��4As�wq�O�UG$�{V_0E��4��tX���l�sQ���ˋ��)�P�[#���\3�5ĸΩ��?�Dޅ,ߧ�����Eb�e�wi��m�\�Ɯ/�w(g0��F�L�R��u��^R=ڋdY��|w�ۯ�!�Sy������%������^">KD�<�%C��=-���5���N7ڗ-�I�U�m{�n?���s��H�qE$��<��=�>d�x5rS6�\X#e�:���o��-D 6�"�-��E8T�z01Y���I4��� D����hi4�-U����� �t��C�sK�s�<���5�d��ߕz�%�P#�5�2�?[CFk�����u>u��ߵ�ǒ�c�(�?�le5��_K���������Xz�����wi�׽d4}
i�s��Y�y=��5,���:c����b��`ɉ�r-�cD��M)Z�<S����֬�s��[�����/H������x�Wi��D��č�ㅙB�H
�I6f?�S�%�F��L�4SK��z�5�X⚖�S�?���Z�<ߗ3]ZWͥ�c<u��8�����%B����@�%"�q�Oq�k}f*�A�5�?�y�q�5����aY"��z������]��g�Q�H��Y��5�����8������g�}}�jB��w)7Rٿ��z�a�%��[|9��F��?�cL)@�	o<��jo&�OD�Jj�>;�w��k�x�~<W����G�LH���9��K����R.����!�V�b���XpU!È�#9'�$	CG�J�+�Q_�w�����2[�]c/{��S�|���ֶ�y=�����S�_ꋷD|��!bED�Ƭ��a��D<ָ�zo�>[C�Kk^��<�wyp-�%8_ڟ%o��ZkS��:�/�-�V�����~���:�f����[D�#�2�jJא�$pfO����H}fDu�ɻ�b�(w���aa4L��՟D��K���m����c��|��c	x8]gM�0E�$�+���1cf�:�H�w�2>�=��/!�5�~�Үq�k\N=f}��֖�Δ��*:�%D�t�Kߗs*�[B�垜=��;K�UG����a�N9~�<��K.��:�8�z��~�1���gk�o�e���<�<�:�ZK|��R����7�ż���m���}/[���x��J�.!�9c�$O�z�q� Q���5E��s�M�p���<�?���w���o�-~S�� q@�2>�l�eq/$��X�m��	���"�~�p�a�F�)�ц����ƞii�}y;K��Zo�"�J��f��+/i�Q�V"k�,��R�K�6ܖ�����6{�\9�p�2 �ߕ��������d�Pr���}��B���g'[����^��o���ӺFo3P�_s�"���垖�]��/�5�=���!��j*�_k��~�U�,�>�<��RD怤���N���U�B�q%��kĨѫ9Πi�3x��G�c�3d�8�zO�y�g����C�!�4X���ku��Iو�!�`ۨkg�� l{<�$�k4Ƃl��A� �a��i��ߧ}���z��pM,����9��΋1(Q�8��C��B�K��}�#�%
���-q�km�٥~���'��a���]}�*m�3����|��Ʊ��eD5'��;��]RF--��y*_PI4�涄����]��{�%�]��5�q�%�������*��>�Dn��k�l鼗�V����%ڹ�W۞��gi��Ο��[�������ѐ�H�+�g}<DĨF]L�|<��S��DL��XP�h���4�I��ږ�\�R_W.��o��@������V���� ^�K��%\kK�>�����l�ܻ>˟�I9y�Q�"~������!�%dR�Ws�O�q}vK�cmG)?�Da�k�\{��k�R�m	)��^��GH�	Ƥ[2�V��A)?+����.���/絴浶vƧw�4k�U={L�x􊋥K=y����l�E(�<�ԽТY�M�S�vVK��-!
�7L�Ζ�Qs�dQ���=:�'.���s��؞�(�/�i�e��.���(�w�*E^{o��!�z���wu�kc�c��-�����5�g�?�USK�jn5�}�W��#K�^�7�[�ZC襊�ky.!�z��\���eMȟ�����k�����z.O���*[ڧ���f���^J+��pZkJ"T3�k8g��Jj��q�}4N�&�a �TOĠ^;B���4L�s�Y��-yh�g
=�89G�Z#��S`��䵢|5ǥX��KS�%�}����w����S\g�쩱K ��]_̿���}�\k��3�;�c� �K�����Vs���f��2"4���_�zY��r�%�Y��e��5\����c���.�h�Lk8���f��fJ�5��=�m)��%j�*��4�#x��u����$�RH�-u�T�v:�:�?�ob�� ;��XLh��"&�c�����w>���BK�
7�
�[rM�9�%��}8����A���k�D��S�/���e~�۬����6��>��a���}+Ϭ���i~�<�5����k��2�X��gKgT��3���F�9��q���޻�3X��w������5�ui�~=%a��.�e}��b���Y��	�_{����1$�_qk�f&�L��[gA��z�,q��\;�|8>�����x�O��@�iQ���������GA0X1X1Qum���'�"���y���Sf��=��7��n�ɼ����{齧��Sk^Z��z��5#�:�s�*/�T���ǯl-��=�]JGk�l��5�T���]B&�|J����d���{liJ�e��Dd����5b�?_����j��|^O��;5	�([���7c�!{{���pn��S�9��FcR���IP�#�EX����J��O��D!x~��0,\�Ŷ�4����AԒ�]�Ɩǖ��un��K\ջ8�5$[r�����B�K�}�-���r���x�8�:˧����K�]&�V#��^������T=��[ת��/r�y?E��{֐~�ğ⶗�_���y���\k�wI����8�:>"�Q�o^���إ!�)�^kg�3�w'�[����j��/�S�٣��)"8��\K)�C���ӷ��`�[�o8�G�-q6���m�v������s��)U_"��F����I:�� �#�m��7���ݨN̼���4X��C���4�<�5�?����s���1��tAc,?D����e[�2X���]N��ı*�q32���* `�}��f���!ֱ���	���3��kh��#�0̟�Y�9@�&�I gL��4j4����q��3��J����k[r�,�AY��C��[s�˚H�k-gi��s-�X�.a�v�,hͤ�Y"L�o_���k�}�Տ^��~+X�_�͟�U�g�{ͨ��s���rM\�18�0�h1M÷��Lt����hEc2�qK�4\�k�q��n���'
Lq�C0�D�;�x6�|���1�X�Z�	B p���h�p��t��� [~��+�en���qR`�8���.�&)/�4)�0n�T'Nn�����5��n�HԈ���K^�RbX���S~��-.�Q_����|�#����u X��Z_��j]v}��GZ\#��K)�>�%��ڙ.ͥ� +�{jO��k�L���Z=n���-[�[�����y��K�����^����U������h�Ϛ������Ĺg��])v���Ƅb܂ɨ�4�U��z���w"�G�n��"%�{�|;�͉$]{qa�C��)�|��B�s�OUr���m-V0�i�N�͕sZ�n��w]��k�P"��<7s�K�.�[��l�zc鹒p�cfϚ��ޟ%��|6G.ͫ�R����˽��|����"���2��ڞ?�����>���x�p�D�F�Kĭ&dO15a(�>���sN���)����*{脘r�ń_B���Td8��IVwr�����T�! 1�$�h�sp�FH?s���g�AE�s{������$q�9�8�9>�}Y$��1Ȋ��E��ԗ�lk�����Nsx:�ߥ����TNg��r���~�6���������,��)�{�jD��<�E�����Ps�庖8��̈́ki��8ߥ����Sp[���6N�\=V��zg�;w=��y��>���Qq湟�.;�z��r3���af��p_	_��fp{�'ߧ2ۯ�>"�S�r*���kn�0��s�DK�VA��B�DM�9�q<j�#gi�v�@�����Y�ӿ��^���R���~v���O�wNϯ��T��م��]��%!�s��F�w!�%�$��9R꾖�v�ת��9�2�!/�a	��G�N=֒�%�Afh�`0�S�U���������k����%��6�lժ�zmke�yX{�&�u9�P 3zkv8�ui�h� ��65ko$�<� ①���`�H�S� !$�F@$Iւ��P�
����!�|�~�1F�			���`��ZN)�SD�`���OSd\�<^�ٯqv�ʋ��K�,q=Oq(Oql�\�b����Z�u��,���8��y,r�8�q����j�ﺕ�_ҙ�!������r����~���A~fI׼Dhʵ<5׵��6���p��iXv'-���c��3ĺ��u��gV�_C���߅$0����a�����t���B`�"����_+N_Ĕ�R����՘����߃3Ĭ��Trޔ�^H>�1q�!*14��Y��e|�8�h��F-�BH�s�@$�Ν� R��H5+��-��b��|Nϟ�K���q�K����q���/9z�	���K�F|p��c�qjK�l�Д�ՆƧ涴�rm�g�Y�[��{���%���ga�{W�ZpV���\�RN�g�4��Y��-q�%��J2�?�U^�R��sK�Y�M�'W�@4��Y%?��h.0�a
�M�F ��UmCy�rM�D����yǼ��pRY?��������=�b��>���#��S
\�M��K@���8�x���c�.ה���]�%d��\��5�欖�1�r6��_C��X���ח�)��G�w�������*����K����]��>������Oq�k�~i�K��]"KU��W6�%8��Qr���g=�rK���\�����}�}�t�5"����,�5����}-�]��%���7ؘ<��<B9���k9�ӥ|Iќ3?��?����:�"��)��b.��߷}4��{����sWx٫w����	�+#JPP ��p�0�#^J��:�0�I4MrN� �Ӷ�|��Xq���$#Au�<�@_#�����\y������9�ZBʏUR��]{���*���B��k�Ps��%/�<�7�����)Pz_����Xs+[�I��x��b��m;;8�ԝל�eo��L���,%���G�V#�\Ĥ.�^#�r=�����J�R�5�,�U�%�%ߩ�1(c�`�97#�&�s,a���S��)�!��ɵ��'��1v���0"�"d�m2�,1j���x8�t���5���bk5���d?�F ㈘ݼ'�����3��s���>*��\�c��8ģ�ξ{�82�f�Ie�\��xf���)�wk5��|����2��}�X�s,����|i��g%�y
	ג��u+�r��J"S���[������[��z�5�����?�3���(��֜�Z?Ks���:�r���^s�K��r�jkDi�k~\�1O~_��T�O����Z�G+K�g5�����1<���^H)-gEIp2�_ߑ����x�>H?N����=Ơy%捖 q {�h���%�?��y@]�֭������U)B�+v�/tQ.l��K��n�+fՇ[s2����-9�X]�sp��꡾(kHH�b�{�w�������/��=w�B*�B
K�ci=�3k���� �%��Sz�5��\{n����Hm�rme[��z��������3>�r�w�T=��Q���{E��9G�]�l��X���f$xO.�)������'OD#��Và��E?x��s>b�M8��1����և�_�Q��uҭ�n�{�yՀ��>��^��T+U!���l���E]BX5�^�k��˰tk\�B�ۻ�Y��6�55H����W�%{���}Ն�����zW[��5b�A�׺t&ks/��>s�u5Nɨ����+k��KJz_I�<�%O��=��/1V�諾��L�<������9�*�꾆���m\6��f��Ѵ���T}&���cL�}d�r'?��Hd�2���#&"�/m3@�g8����^�%n�\9n�a�g˪��k[B.K,��M-�jD\r��g~�]�$����R[C�e��:j�Z����H�tn�g����bP�$�N��V����>R�!y�})��Y��2����S��R�k��lm����B�˴!Ɩ�Cd$0�`��Oo�ġo�>lb �g��|�$h��rX�\;$Ƅ�(�9��|���S+?	t�w��_��q~%��!��zG��(����y_n7�����F֥>�"B�{K����)Ķ�����z-K����[���u-���=��g��t�\�G��w��.��f��Xۧw��S���3�YiK0�v��c|�$kd������G�s�)���k?�h�c+4|���QCn��,��Ns1F�4������U�
0L��>��}I��ሠ�#���	1LĨR����"j���8	(.G�7j�$��<α^�w�]�v�V#����*R����v���ɟ-�P��S��ߏ��Q^������אm}���|oI���Yf͜	����<[�����]��5¾F�K.�)�\�����ಞs�ͯ�c��/�a	�K0��,�:ߧ�5�Y"��y���	�dU��s�ok-A��h��>L�:K\��_i��=$O;�5���)r�)��}�QC���8��K�T�q���nKW9��gk-�����"rf�(�^��2��7�׷t9O��zN�u���|�2	�	�j"UreO!�z]5�)�_��g������[e����1K�r�O�S�s~f)�mY-ͩܫ������ޭ1+KH�<��g׈�S0�D�J�w��Ҟ,��$cq8œd��iE�[j9�Ŗ�+r�V�����L<*��!��\��5��F�; fK-�tA���>&c0fC4����ǅ���� �1Ŗ�o�xF�����i�r�G�tDoi'�n.T�;��@�u4��Ghϔ��0g��ri����͒�sɽրc<3�ր�}��1̄�aN��R����הו�i���s��=�|�j�Zε&�e���Qs��u��҂�y���J��g��/���1m����0��]α\�R��ؒ�P^�<ϼ?K9V�`����#w�T��d�B3S$��b=��a~�\c��_��IP�F�\{�S���wy��o��7���!�ό�D�\Y�̋F���7��JR�߇i�5��̈́�o1�%�	S��������M�蚎��X�x��=�4c�B�b���=���I��E#f�1���q�adD�#��k��O:��"��ÿ���W<S�`�{��_��4=�3~�y��K���d�bg`^�ϧ�~:��Z�R./�RI�r~��$(���̘���Y.>kβ�l���9ĥ9��.��n�S�E��y�g�{��_�jXYk����<�j8���<1e�5�[�r^9"�vb8�[/;�k��{KRN��3U�W]Oxi�\���r�z�����ZK�Z�xJ{�ML\<�l*��������8=c���9��*��w��1N���h�����!�)���^,�E�%�~
oā��d�=�hȷ5'A�~N|@nٛh]�XW��˿�g�"���S͈8�a�/Z����\��<��,5��ڡ��U_#2k?���Sѧ�g-I,��D��_�����Sv�����j�yW�������K�w����T?���au	������S�JM��;R>[?�FxJx_b�`/�f7�t��'D.��h�!��_�'1��Er�%
��5Bt���1#����#��-�SϹ�P�Ч����9����.�ǈtِTJi������ȵV,�y���{��^C�5�)�P.�/�W�Q́�}לe���굮!�5���`�>�"u_������%��~wi5�|���s����[C�Ƙ�S\گw�/r*�X;7,!��y�k_��%\�W��S�]��$!�݋z�l���Ҧ��2�Z����Sm�.>���g#���s�:��_��_~��т�t�c�t�Z�J3���� ��x2l  h�|3�'Eƹ�?�Ƹ�&4���K)¹>�l%�,m|�ֈCy�5�[ڗ����N�$k����9�r^p�4�֙��'��EYSa�k�=r��D@ʟO�Eά��SD�}�\C(k�/�����e��pi�K���ݵ��	O��ދ:����U�ݝ5�`��έ��|7����\�R2��=x�,$@�!#X�8��[�6)c��gB !x�ƀ���O�'�~��9�b.1q�"3,����>����Z!�p����g��U#�O���{�YK 0�#f�9C�g}d��`�:�%���~.����*�5�qm�����-q@% ���~�F�O�q�3.�}�:�Z9�����XB<��k�di��r�5������ ��]���C�����v>��['�+��Ҟ��Uz���˿kFk��ȭ��L����1(u��ΜK��9����tIyĒ��I�:��Yv������}��O8N�T�����w��M@C�ņ	���n�(�#�WOIUf�����'�|�+#Ɯ����F��	����T0����Œ�b�#.���������S�.��>�^_���%m}A��|kU��k�m	I����cן��a���a=5��-�ڜ��_gIZy�}Y�n� �?e���$�w18�xk�A�_�����sϬ�|���S*�z?ט���bپB� 1�A�Y�.��s�UZK�X",�18�HD=-�@�k-��Q��R���N��hz(g��/m�$�,�<��6+�����\|zZ�W�W%2?�����"�u;�)iT����K.�|�O�V�ٔ�\�OG��?kk��,�����=������KȸF��|�xj�D(���.���G�AU�����9���k#s�lV�-�]��~�u�]g\����*�%3!��K��.�^v��ʛs5gN�.&��O<!ZӞ�8�Tя�j�{�5�H��J��U�5�P��K�q��81!`74��K�����*4"���i�� f"�=�?`c���V9T�\�pTC����V�S`��q���XhZK�3M�ړ���'�9�_zN�Dl��
j	�J�e�4�s�5�\��-��i��^Ku�T��ө�Ҁ\�vqK�%N,�	,U���>�aTs�����W>����iμ��2��w3W9��ꭞk	35l��z
�<����k�j���0��2�{>�wq�5�cp��'#�)ϣD���K�W�	Nug�z*��/ם[��ړ���%�ok�[�Q�����S��#���Gi���%�H��M��[�T��m[&�H]�;)B���C��+1 ɦf�J~�LS 6�F�|�9&�X���=-�0��Ɉkʀ��/�.�L�Q�N<ҧ�}�dr[�p�5���{�xˊ�^�[��>��}{�i�iP(F�c�|F�C��3&�!j�KP�$���h�1�/~p�`��<0@$�����ݷ��|��w��ګ����>�"}���>��9���Uk}תU�hq)�<%��$wuڼ�y$~��eTF�U��1�BF2s>�mW";ɼ�d�u��<�,���~���nU��x]H[�$�&?pE�7�I�ۣ�Փo���-��4i>��x]%���O�+2gС�iX�R�	�'�ȸw���ϸ��g�ֈ0A���x�A���b���zYX�6�6YDt!8i/S����L[g���bǜEj`kPhFA#B�&]��S����/����kePF�_+���h�mF�S,&~��P�6����&�ס$��1ƣq>���YE���=lS��$�롉-��Ѳ>UyK�!��D�2��:H�@	Qˤ�;$�O�9ྴ�J�ȺI��epf�U�":�̹$u���*fɯq��U�lR�T��W������G��K)�{��� �:B�\��=��<8��:;��0&F�$n]�w���`��Y�E�ac�Rc0J^��"m�M�Z�={0 b*7P�4,$����&�:c����G���lJ��3tYvH�b~��J����즫w��O�ߗw�D�b���*��U1��;�:�k��g&�W2L`hB�P�L�7/���s�irf�J(?Y6GΔ�N]�尼B�wR�V	^�$�"�,���|?�\h�$����h;���l]���9�s(�����v�1n�*ʥ2(�~��_��S������P0��T�� E���Psb�>Qnu��Ո���1m
/O�ġ|3�:5H#Ks�E� �#'���r����h��4`�����s�Q��Ǥd=&!$���]�e\
!�*fV5���$��|7��Cm��[U�(ߕ���8���sFϑ�$�*O
TY���]V�����f���֡[v���ݑ7#̹V�5�+4��y[5�Bɯ�آ��YPX����@gw[��*7Y��s�i�TGά	5`T�_h ��w&��ºC�?o���r�e�?�����ֺN(�Z J4��H�$8�'!�=ÿ�P�d�����Q�$�YUy]�i2w=4�Bm��cҒ�I�ϑi�������']��G�k�Z��_���Pv�(�:�a�I���$��P;�"��S
��
�*Wg.XB��'��{���I�&�������\��f�ƲL��ضy�����	��$�� �Xh$��0y
U�n`"X㤝�5���&�:�N\�k��>��.fL�~4�T����d���������ö�q���QR�l_ʼ6� �{T���3��U1�q�������������7�2)�\�F��#�JU��<BB�{��I�\U������tq�}-����v.k��%Pb����h��o��]�o�p�eQ{�ÅN���Y��|��8�P�&����
��)�
q�[�����jX�\�0U�[Z���eH:��ygK�0pGWR݈��*'ODL��(�1���d��z��$����$���{����̪|�����Z(�qI�J!J�z6��e>�r�y�⼜*!B�,ːeYiA1��ƍCH@Q"�i*�=�,AU�3!�%��d�U��Z"�*N���%IcrxR��%4�\��n�ҌY�5X��[.��3��j5�%����Rj�s�̀���������,Z�:�� }��&+��T��Z^6��s} �p�Jtd��.���`k��E��`m�)R��#h�^��v���6F�h�c:i���б12��W���D��P*-�Uaf%�U���F�9?�D���W["�a�a���-Q1M�<eX9IJ���U�����>/�O:��Hͥ����
��:�g��m�V+�_�m�{/��Zc0��h ˜�$	��~�q��*p�w�!�LC���'�2��B)U�oh��la/7�޸R�x�=��8���Q�BtH��]
���e�yM.��~�
J�P����}�b��ڋ87�:F7ɐC�^�#B��*D��,ˑ"�6��"�'�á�<jC�	t6��@7 4�O�hF�Eg�s�E=�C�)��ذ?��M1f	l�1B��'m�����Z[#QZ�T���	5�`#Z��<RSJ!.��i�� �܎�a?�WFr�D/QX��"	[�/��	H�brU���=N��m�L�_��a\>!�$*_-��������h�Z��i����Ś� ���Ҋ]�Μ�I� 8�ߏb�{�=�ʓ��_�J��D�<?ʓ��Ծy��ʪ��'�~R��^U�>1y)�dY����1��</�Y��|�h>�g��G���xZ-D�����4�~���.���I(��` �J�"ٹ@HC�҅���İ�Jx���-"{:�}��o��B��Va�gV��I���V	
N$2ɅPIJUO��s���M��b�}���̒����⩍!�E����l6������$�}�n���v��E�qއT���j������	哺O�"1)~-d[�B�J��\>�h5���
0�������P���k��ǁ	h�6[>��,��px1�O�!;�z*57Y�~}�Lζ���شULT�!�U�<Kt�=)�i�^�7ҟ�'m��&�H_C�J���-Z	�uIs����!;�x�B@��='�~(���'g�2�8�*_�&�����NB��
ͅ�^�1����K�- ��}cc�zq#�2�j5=z��P�	���%�kʄ7���Cm�D���y�l6������K�S�ϸ��}�bv2��|�F���W�t�Y�jo?/?X�<Jr���3��4�J�W���3��;��8�8����G d~�������d��L�"64܊xq�U���y����"L$�T y��o�58M�*%��%�!���zF����bD���6d��C2r9Qy����
��q�/�-�	'I���i ���j��_ch4�Ij�d|����W��z������y�C4��*�)�I� g��9z&dc�ɸ91is�?.����q�'�]PB�|�D�R+M!�h�����;]K��y�X����* ƶ�?�*������@�^k���]�r�/�(���8�Z�R�-�G���I3�AGБg�j�(���j�Dk���w�0�&?6�9�ߛ�DT�Ld�r��+S��p�z�Onz���b��i��~��8�p���{���:�mۆ�����ɏ�[I�	�*T?�FN��Ly�z=���x!���F DU��C����<e[B�$4���wǡs��SH����>�$`��F��>�#BD�;+�f�/��y��m��2�C�>�2�I4q_�oΪF���bkm�t(����	j�N�� ��$��5�"U,�pG��Q��
U�י��{p��T��LD%��T�M��9�yȉ�QM������⮦��-�4�/�(���z�V��?�.��2|�_D����[�^G��28*�e�WQ=�7G}���5B��V��{/>�����o�&��XJ�����aR�})O�
���j'�g�T���O��~��<I�v2U�ID�ي6B�\�Ӱ������TJ!�3���͐�)�<�}eea�#:CX+s���oll�����~�����p�{�l�} @�A�<(�!�ZBTJ�ܛB�*�0�=�B4<q,����Ⱥl��8;�,��BT!;�d�|Y�G��<ϱo�>������ǡ�����h�^�������	�BhR�/���;/���������x׻ޅo|�h6��C�3d>RP���P��_|�]����	dJ�>�O���
8p3^U��$=��6t�3v9_���Gx��>�eUi8��Zﳶ0`�����N[f�q(o8HI�@G��J)�Z�K�Z9B���6�(�����`0@�:��
G�\S'��J��)Tq�YE0Y�q�EU�'ӀK�	�YKB&�(Ib��@�-x�a���u��u� ^@�"'#�x��ȍg!���>%w���u��udY�V�c\��z��>��X[[s6�z���������z�/��8��D���̌��I�m���*�I�^G������Zcyyg�u����_طoVWW���P�Ր$��P��/��/=C�F$��k|�Ս�Af'��@cbz�/�Y*�����≗O4��2���5NR���B��|�y�k/ѱRʏ�c�$P��ځ�c0�����ˇ%Yk�U��3)�`p�O��K��ȕAԈ��^ck����5f�����*��rn�����Q"@c��wH��)n1����s�ZmKL��;u(lO����������Bτ���Q��'V��� �:g�9U!�PeB}��}I�:�x������g�4Q����}�kq�i���~0 `vvKKK�����o��&�q̉3��tQiS�Qw�]�A�뿸��;vx&�gڜ���P�d���	1@9ޜ��v �x�qO/�\Ќ�q��o��Cm��K�����,�ܾ�Z!���P�N�Mńa�eȊ�\�Ú�R
J!e��c��_�����״�a����9���j}��*��X�ڟRO�z�(�;M^#�bh��Y[F�.�lS�1�q�HU�A�&��q��8�?�!�|���B��$�(�we���n����)���Ak�v��v����t�]�x�x�ހ��ؾ};���p��!���baa������a���Gи��d�ɶ�q�=Qa}}�f��z+����� �OS
Y�D�Ϥi,ԯ�������I��ƸP��/=�1�M�������5����u%�3������8�o*�}�M6 r� r(=A�0���Ï.�l*�^@��s���i�X3�-ݑ�Ty˸�e�j� ~�2��k�X�$j&킂(�A,ɟ����"xW�0����dpϨ�{��;��U��扪z��?�d{C(/�*ǵ�L<����򗿌[n���K��n�g�q�mۆ��3��g>� �c��x㍸뮻�={��)�kWyj����:�q�u�h=MS����VWWq���]�z����=�Q2)��"]lC}=N���xiR	��<��D��*��?47���8��@jV�L~�����ma���Мi:K7���ʋ1�cGJ��1�1@sC� #�ڱL[��i��b�*����$*Y��Š�P{�W�S4,i�/��.V?#$�}��wƣa�^��]
�P�����OB�U�_-�ʶT���ȍ�C��f�I�V�&�[o�_���p�u�������o}?����7�	���7p�UW���~7�,�7܀w��8p� �(B���$�c�����t��?Uh���֩��=�܃o�������N^Dr�{���"9&�.!F�?��2!���H�ޝ�BڝԘB(�
�s�9�R��פ�4ls��'����z����� �\]��( Gi�k�q�Z$\E_�C�wη5�m3�f��R�P��<2J� c)�t��l�QJ��3%]a�_�dB�y��a��͖'��E�q�%^Wɴxy��FM �o%���&�Y%��<���VVV�ԧ>^x!v�څs�9�������{��^�۷KKKx���Z��.� �w��Ν;1ܢ>[��ѼNR�R��-qB2B��V�nsssXYY��?�y<���.3S^Ӓ������O�2gq�+�k��\&�c(Q����PY�>Rp��q���]����P:���S%x�S�"�HA�" ]�:����8Fn#]����zS�%�b��1jA��p����w*u1��;��^���E@#e���X�j�a��Z�E4k���7�s�p����uڄ�C3�o�)�I)�*7DL2?�C�b�|!MN�O����-�R����EZ�F�!"�Q�x�e�t����Z�;v`Ϟ=H�sssh6����q��ף�h��x�<�L�}��x��=�AX__�`0@��DE�}�X��Lbj�^�H*ǈ����wߍ?��x��ކm۶���R��B`A2)J�)��BjY0Ⱥ��l�A��{�~��?,H�����?��SU��Uǅ��
VIG�<�-��N�TL�F�X����v|��Y0ls�����@�[f�!��
�F%"	Ha�Ѱ�w�IA�R�OHU([eU^U�V�P9t�
��ߌ9�������k2���8�J�	Qܚ$I��v����4M�����ۿ���í�ފ,˰���v��~����%,--!MSLOOCk��V+�
B�`�!'�o���Z-��u�ڵ?���O|W_}u�}���6��:U�)�:������r�	O!аY�/�$�.��!�O\�yF���z�V�����@�l;�n���R8m�oȏ#}�w���o����/iː~R[@/���S�`q��z?A��b�s� >	@����Al#�����燑�M�"G�C���*;�HՐ'M(�Q����5�(�A���0�V1P�P�Hc�n߫O��q��'W��D��������h��l�[���(���RYI�Q����rn��d�-�G ���nN����|��=!!l�R�L�OL.D���E'ANR=zy�C���������ߏ��9Xt�$>�yƐ9�&dh���7����]����i�&v�5l���h���Y�#��i����c�Z�*���`���۫���Z����1�Z��<ҏƒ3(Zt����D�p��M:P��|�?L���H�4�Qd��)�A}Wd�f"��Bd�l�"��I���a���ch(�a�g)�JA7"�m
c�0P6�z�h���Ȓ*I�(�v��n��NC��Zo�R@}f��H5 [C�.��a��@m��6�:C��`�`�/i��0���v��v���"U��_cL1�p�%����aHB�M2��	1�qH�_�τ�Yh1��U�q�׫��\�QuI�BͲ��C!Ƨ�F���M7݄���m��O~�N8�^y���8���N�?�o�3\��> ��H���&��N�z�x�+_�_��_�?^O�c3�'�MZ��u�y��i�!̓Ө�\i�Ue�N���&vt��D���e��� �'�Z����'ǀ'�"�i:�� �2`0�*��d���?u�����黅���z��7���������*�>$�#]D�0�c-"��D��3<I� ��󕓎�~��>v\�HI��_Y�P��C�-���E��T	�P�yQ>����#G����^�7���˸~��J�/��CϒY'�2��}����?�)>���ꫯF�#�=!-/��#4n���U��5i�u��ו�w�\��u�u���P�����	FNK�[+X1���&�\/k\���-Rfy����Cko��s]�7�5�_�5
.^رK[��Kk,����r�tI�Ȅ3E$ng��Ƹ���Y
�$����!�L^1�/2�3�/iR�e�6��d�!�����q�\X��H�	�oll�	Ox���cvv�n�Vy������6|����-Ԏ*������6�:�S��8F��
z���t(Q-�g>V��e�B�%�Hh����Ȑ�Oz���\�����Z[
�Ǔ�=�,@[m�^YH�[ܕ�R�9�� �s�<"=49��%~��*����ts ��f�3�^��$�!j��[ȣ".E�t�����Q&����6�?X�~��j�A�yk�)F��X9r��I��&S��Jց����B*�$$�0����S��Z]�]��P^A��*�G�4w�؁����C�b:�Y�c��]���@���V� 8��&VWW�k�.��-o�`0@��E�e~�I�qS���4UI2S�w��>∼���XH��M����3��VD�y=i݁������S��G5�*�ܙ�qd�P�z[X[�s���+����X��@�����%�Ě�Hj	`���Qѭ��cDQ�
ք����-�V�Cf2h+G
�D�Dk��Vb�%� P�R�E0ef)�VU���è���̂_�b��a�|7�Ы�䶌���?�)�� ₢V�y;��W�\��~uu՛r�,�EDDi:�B��h@��2E�5bJd����f�	 ��/����!����4�TцԗRK#�+�
%�F��׍�Q�x��ZՖ*�&�ͬ;�Ik@�CZ26�������~EL�M[�]��2�P��(��RH?�ct:Õyc�v��V�!Ea�W�ې뤧!����p�� N%be��������-[hRʕÈ.7��D�|Gi�������%c�Z�����������7�~�m�z�0�~�����:�ŉ��)E">i��,����}+���n��(��n����
c:��_p&#��)'tH��s�L/����zO���n��ӕ��LH����!D!�^^�3f����N�5E	��p<C��cH�(�T  ��z�`���Y$q��j�e`M�F�CI����"�رc�[��[�����8�F
3��	�z|kE�Q�RC�p��9���v�4��Tn�F%A&�UUi��b���I����(!�*[�*��/�'����qZ�d<����&���肻R[�Q�WʝHEh0�|�yra�j7ch�%����������KKK�}tcc�k.��9���y\�*�VՏ!t�]%��"��3��'yqaL`Cҭ�;�&�� ���Uu��I�s�M^*�}�>�����E��1�0�N���Iı�H,�)b�ZK��Aw,Ӗ2���vd.�B`5�}49Z�؅�!&RĿ7�Ǐ���(L�#��m����6�H�z˙ �ۦvv�Ԥ%���Dn�R;C�c���1P���Q������`��/�4�;�l���4P� � $�x��������4�y]�^�P���rQV
�$I�k��;���ݫ���,����tE,1���d��{��x�|ޟ�dB��Z�t��L�6�I�B��-dKm�*ޯ!K�gtr-D�%������r����@�׃���*��@NN'F��:��#�A�"� "(3p@�*h#)��~��T��@Ai�(�V	�jp6#@�:`�# �.�&� ��`���9,z� F���ϓ����z=���/�)]^�O���lZI�B�m�=CK�Pgi�B,&��;�)�P�a��(*�C�E�"z�n�U���%򕌷�ݡ�!�#���OUm�l}d��I,'jU�B2U}�W2�*��l��߲�r�$�TJ�ϸ(�����B��~����V��
��lk��B�Ɵ��7��y���W=#�o�,.W�O~�Us��R��ba���eYU/N�C�P�@�vԼHut�`�B������zҖ1�4M��֪"]�#�`5r(����A
k��5f�;�yA**l�F�S���"W��bal�E`t��ym�G�Bn��2�&��زr��|CB��G^7�Cu��Л,��y�:�&G|!�jYF�Y_`hJچ� "�����R��j�>���%��|�4~��d���wH���~�8��3nބ �!m ԗRH�6s�)���@�Ӭ�2���4@����W {W�<ϡU�(zdE�F�kP��T@A��䰆��W���EDMh�j�;QKGЪ��Yg�HD������s�e�PV�*�r'	�l`�BLDk��6Q��z/PT�˛��E!e�3��C�UDU�r酞 P^�*a3���lOCMdٮ*Dj70��PNj�(�z�U�H��P��,7�֍�P;��8$�˩�U�B���4)��H�J L�3U�U�^.�g�����B`0$�H�PJ��,�����&g��Mh��b�ҙ���/^G���,�x��B+[�e��sJ9�H[�Ѹ�942(FQqcb M�d���
�78:��$	rK�.XP1�p*������D�(�Jb��x��I0Ĕ����ڡ�]�?�UMV�l�0���}I�b%��*W��ǒ�$�'�2��,�����4�4���ER��t��|�����|F�y�G6�*�,�]U^w�悛��}��y��T�irS�1&xz���6�;]OAi�C)�8�� G��*Bn��V9P�Ӿ$'�#hP}��!w���,���J���F�mC싟'm��,k��˔b.��0OÉU�q7�(`���-��z����PYU����ơ��wLU���u����*�u_����*��x�jS����U�j�6$�)�,������SY�P�)Y�|>x�U>����[	NBm7n����S���m�2��r��P:ra��qx��Q�a����|2��ga��g�~D ����X�-5��'�	�6ޤi�F��ᛂ�G��R�qQ-���m�
�f��	ED,aft��&u�#�ɈX���TV�pC̐�5�X�s9��j��#�'8�!ѻ��l(�П4�q'��{���S�&��yݹ�G��;ңa�ǵ7��q�#{>�>��Q>'˓��y^�L!z�����h���0uV�!�qB"�@������-��)2idP�<�(��͠l��Ӎ`�.���@'F�N���'��%��~�-��1j�!�X�m��.z��(A='l"x��92$A#U�yU1�a����*�;	U�wC��:r�y�c�rR���K��
�Ф�H��]�7Uυ��*�@ޟT�\�� ����+�����)��)ne=�h@j��Cu������q�eY�t�}�I~?TN�/B��$�
�
#p�t��� ��C<&�X�K⁑��uj���O�2���#�}���X��\�`u�S�`"U�� 4���9���L�&����@�qhm\q�F��1X�R
���<AE����߯5��6���ܠ�j�Ƹ�m����E�!t���1��_�D�ôn�w�Uq�G<�>��Uʰ��nHN�҅�|��}R�����Z���O��vhz������+��Tjg6��,�ny����6�vk�?��v��.0u_�5�,�a�ܭ)��D
TW��R�V�m����%�͙8g�t� ��:FD�����[k�bs�"���ǧ*�K��F��1C��Z4j5�B��Ӻ�񹰹�{!�[�1ႰjM�m3(������ ��O�3�}���l�]�����*�1ȣ)�+<2H���(Bf�����I����Ɂn��z�X#�t\<oz�@G��Ы��:���As�j��@���F|�1l�w�t�S��V��e��J�������L�*&M��R�i ���8�>Φ��v�z�6�{�����z��I�F�`t�׋+��I�x9���[��'<1M�7aR����)`�l�~b�$X�f�Qi�N��F^G)Cc@�j�%S�����ۧ��4'6��h�'ȼe�{TW~��_.���;7p:����6�.�_xd?:a<l��ί?�c(S,BS�b׮R


Q��������њ����z����y����}_��G��aD��� D4D�4 !�.ݣ$=9��j��6��O��Z�W�_ MRN�U]2�7�\��8�F#$�z��'p>�8
���+�H�	я�o��P��o��Io+>�r��}NO!�I�A
#)�B�oҘ{�"�K������sq̚I�>����;�-�H�}hބ���`�f`���Q��]ynEN)@��>�&��" $�=��U��/��漊�V�9�_�e���)��&A���~��#�O�K��:u8��B6n>�$S	�'d���Q�l�"f��"/'D��>�1��T�&+ˑ(_��BL�'n�QlLy]�}$Z1|*�L'�v+����$I�(#p��I���D�a\YG.�����tQE���1Ĉ�r&�It��G��q�
U�C���G�Q�_
x2-JA�ː�����;4�<T^�E[������(�<�����֯�s��zӖz�h]�d�/�>%��+��;�~]�N�l\�JY�������D����&}�I��K5\����ja�z�gBȰ���,X�.�D,4	CL>$t�o�_.��@$�#5��B�!\�ҳU�W2Ψ�f���J�����#f��q�%���
ٳC¹J�ɾG'�����(�����P�� �|^έqN��˸� ˚�G���;bܣ�)��yc3���F9_�A�f�`�aI�Y�ѳ+3�&M]) �,tT(ǒ�S�r�M9Х��C�Oxk�'8�3�RL�*bm��`�M����K��t\՗$4��!��������1Z�Q�ɟ���1�C��A�z�@m䙕�y�pxަ�	<�%�d��z�^)t�\L�<dy?q5�%�M�/�>.Q�r���8�\ER �$�?B�L2k��	��*�R
�I���<�H����iDk��3E��`;�r�3}���!�fc Cq����ّ�Q��Q[�1l��-��Q�r�O��N4s�k*����}["�*�x���D�I�w�$��H�-�U���#"����?]�y��Cu��r�,7�p�%/��I�����H�W��Q���,dB�K�\9����L��(�� �_TN��G����ӤB����#b���)�7��r�%����!�W��y�Zk��=YϪvR�$p	�d�r.W#�����������@#�-�5Lf���-�ס����Y����Q%^�+V�jg�ϓ�Sm��|�nR=�KL_)�]�Ei���4�	�
/Ix�P$#�~9qKd�	Q��U1�A��=ʯ�]<O)8S��vjG����AJAF�~�_�2ȥ�����1��z��#��.�~����� `}}����^���Ylll���z�z�8��Z��(�0J�@��'g����^h�#T'y��~��k�">�G~n��IS�y#�������*"�e�f�39���U�=^��e0��1����@���)����(�
���47�oD�Uڲ�YNE�9�~�mֿ32�^Z@��q|t��LLqR��aa�f������)g<�W�>$��1#_>_�������ʅg�6Nm%��G�(�GD*��������.���/ǿ�˿�ӟ�4.��R=z�V���)bN333���7�����7�j54(��>P�}c���������~�����^��;��E���;��V�����ꫯƽ�ދf����]YY��wމZ��#G�஻�B�^�ѣG����	�Ç��n�]�I����$A�$� �4u;ʩ�~�#=�B�k��`D��ȑ�I�4�h|���4���Mf��化Dz�Ӱ�[\� ��~�zѾ��P�5ʇ��f���`��k�qq��d�~�5�v�]�$�8�C)hU+�Ϡ��G��``����sI�ᱡ4��*mӧTB��sR
1\���w��r�$�@���U!��G�wC�g����u��PB��*�=�BB�ׇY�ajj
��qꩧb~~{��A�Ղ1�v�O�,˰���f����E|����=�܃��Yofi4X^^��֣�f��O~����' C����^__G�VC�^ǝwމ�.�_���n��1����}�~�����_~9>�ছn�k_�Z|�����.��2|�����:������0��������E>��O�/��/��9v�؁f��i��F���w�9E�!�WT�� �8����I"�t��	ѠLr^WՅ	�x[����C�$8��+����3�ɛ�s��� H$��4-6o����i��;<�0��v�T��
��P���E�
���NR΋�#�c���ߜ�C�j���n���B�v!��z����"��y9��8�����޽{��=���ǳ��,�z=�z=t�]�{��t:���B���`0���"�=�\�����u�l�1���$I��v�1^��ס���h���`ZQ�~x�C��@��#=�R8�������v�������$	��ۇm۶avv�w:����177��'}�(¡C��w�^��������4�n��&���?�/��/cvv��˘��B�����:�ͦ��XK0C��U�i:�aHڒڭDʜ���PB����$����z�~��4�~q\�Ø�*w๊������
�-t�(0�G�q\h¶��d.@k��Ξ���d���x
��_����1L�)L�p@
oFz��YA1Il�-m_�	Fv}k�qؕR�є%al� �}��8�̯I��-T�B��tW�s\�Ue������v��d���G?�k���Ї�o�>lllફ���f<����s�����ySH������1x�[ߊ��E��կ����y|��_��������>~�WKKK8|��7�XkQ���l6aLq�&Ckqc����t:>�B���/��/�?���xի^�n���۷���=�8F����_�5fgg�׼�v���xӛބݻw#�s�ʯ�
�����N@�����������,W����H��Ǒ/r�q�x�5�tC�I���ns�\��.������_�����Z)�Eҷ0t-�"([����g}�#;n����9<E{���$�md*L6���l�vp�Җ�wxA�%���/%C�|V�#f��7��<��chC�yn]\kKg��l�-����&2)>�&��Um�)��V!��"�P���7I�ձ�M�$VNp�<�D�w�y����}t:�~���b���8���k�.�ڵ�����:�,���:VVV��/��2!MS:tkkk���h4�Z�j�������u�x�l6E<�������W���<;;�#G��� >��`jj
�NG����Z����q���c۶mXZZ��'��v��~��s�9��~:���/�+�@��XXX����ݮG�������<B�g3c�|mV
}.l��e�<1���s�~����ܹn1�Z�\i(E�8�A�re�iU����9&��-6�I)@��ZkK&_�����:��y�cG�"Ibᔘ���e�gX�tJ�*dZ��D@!��Z��8�\%�%����ϸ2����B�@U�-��.���E���?ƃ� :t�w���_�Ç�����q��'caa�/������h��/9�9���o�8����G?�뮻 8���*j��"�����d���Ʈ]��7�	;w�R
����Zc׮]xֳ��SN9���^Ȭ��#�"�j5,//��z����e�ޥ�%���c0`ii	Qaffkkk>����B����-�I��V�&2b>2o9��1	#��|��i1!�}hnao%.�B�"�j���HТU9o.��1��Xȍ��0����T��}Y̆ﴠуs�o�O[ȝ���w�݋��9��)�k �_w=�\^J�$}$:��uӮB>!T>����J���zU'Ġ���y��0��t}db�[����j��[��������Q��077�=X��_�]tn��&l۶ͷwzz۷o��?�y��Ŀ�˿ �c�����������}h�ۨ�j��jH������g>��/���r������h4`�E���m�݆������`ccJ)���x�"��~ �����h4�����{���/~1�:�,<x����a�CL*��p7`�����F.�R�rA��yf��B4)�\�{�Z�8-���Mc�.�:4���Y��HS�3�W,"�kWa��PFx�Z.x�	1ߦҖ3})1K0u����a��wr�?0Y��J��������8M#D��R�W�/�c2n2ݗre�U�e�V���:N:�$����S�������#G���SO�+^�
�z꩸��{�M~cckkkضm�>�l�ٳ����o�>�ݻכN�,C��+	���E�����h����IG��>�)�x�h����zؾ};����g�g��'>�z��}�%Z�v�AD�666�{�n����;.��2|�������X^^F�Vq���J D����1�;����L37~�&:NhQ�^2����]��M
YVU?�{$����s�K�v0�= %Z`k�%�h��<2�83��M��;�^Aj�4���0�ϐ�}��з=�S�������Ѐ[�^G��L�5�ش���a� ���y�c�ȑ��m�ݤJQ�^�)D��wM�>wa���dБBf3?`@9�
 ����_��RMuj:=G�����	�zU	�*$F��ǭ��O�I;���Byp§��0��'1
�`��o�����,n�я�/_����g�35��G����r�:����F�ф�@'�?�=;w�Į]�������p�����xj��W�9'��#��q�8���q뭷 fgg�p8��'�'XXX����R8p� p�e��`kq���P���5�Yqu����i�D@\s��y����*NܻO���bϞ=XZZ�}��v��j�޻�#��<�����z �t���p^�H�`F6ϡP��WB�UC�e��10l�M��J:	!g��1� ר��*���5z��ט�s��Ɔ��Am5tb��֐E5�QF'�&�R�)��0���Ql��V�)Ԓ)DQ��(X�bD1'�9	0{`�^�����bh;�,t�C_i�I�ـ�3��c�#wː>1�*�w&!T�O�I�+1�$U�\�#�$���T�&����Ջߧ�廡����0�wx����yg���q�ji�����t:��w�u���z��g?��c�����n�	���W�?�v�܉��5��� It:��?�3^�җ��_�2���6>�?��?����6�Z-�i���54�M�����+�Ļ��.|�;����|�[�B���6����+�����=�_`۶mX[[÷��-�q�h6�����<??��Ti�k��öm�p�g`vv�z����}	i�����N��㴀�r�]N!$=inH-P��U��f�$+ߗ��5����X�&De�]�I��z����8�m@8���M[����Υ�5�u
�M[H�qUӀ�ar�� �;ir�</�|���C9�of0&��9�v�Y�D�Ԧqi3@�!�ݤ�I�K� E�U�l;��}3�s�W�����������x�k_���;kkk~����⑏|$��ַ�SNA�eXXX���:��(��g��g<�x����?��Q�z�Gx�f��V����idY���yo�'��^�cnn���S��gY��`�o��^{-fgP�4bX��榧�b}y	�V���kh�d�.:�&p�n\w�5x�ů�w��]dY���/�Rh6��Ijg�h.4�U48�69��i��LxRY��r���B��^�;Tn�[P���R�6GnH�0̈�gl����$	j��U��:1mʝR�&�lJ w,Җ{��P�����E�Ӏ J��u�;�;̳j�L��U�p4>*�X}*�$�/�N�9����'��ĭ����s/�I���޶m�<Ǉ?�a<x�����Y�9������+++��G>�$I�<W^y%Y��<�98�sp��a,..��l"�c<��χ���~;�������OG�^�u�]�}����x��E���M]�_=��6N?�t��E/�����6��ױ����;_|1v��齂v�؁��E�i�N����U��}��w��v�8묳p�%���SNA����|ї��^�_5� JQ29=��Bt0I}�c��O��#ϩ��'��ܤSUB����i�v�����1�����P/��_��P㥲���@� ��|��%P��i���u.���5s�� Y���.�N' T��]�j!�

ں�h��"ka�N6m��2b�m�w�<l�WO �`�L���Aώ� ��B�qʑ�T�*d)5#~}��Q�W��k���`�3�Z�����Sk�a�O��=�������'>�I�����k��W���o�E���uqq�F7�x#.��|���ſ���㵯}-�����N@E������[oū_�j\}��XZZ��������f����%�~�阞�Ƈ>�A����A���?��?�����v|�ӟ�{��.�{�~|���_��_�Ѩ�_�<^��K05�^��s�9޻��-
�2w��_���Ui�r�i�C�Hz�fJy���,�4�Bt,M�R�PQ��^��&K���"��5%!S��0���nOE������?Yw����'�;��7�T�u�N(>����1��V���>AŒ�X���o9 Yp���L<T.P�P��$ts(�ϼN�z��|&TG�w�?4�!���f�E�$8|�0~�~�[&�~q�v�����:�<��^�2(�6I��E/���:��永�XZ�m6�����;����p��կ���0�j5����.�<�L�q��>T���9�ʯ�
v�܉F���>��سg�Rޥ��eY�pR_�y�СCX^^F��ŭ�ފ�;Y���o����}=z�m�Z^AE����`0@��E�� t��ҮN)����&&�5)ܫ ����ʩ�	z(ϓI_�?Y}K'YfU��/�n�A���rZCT��Ȕ�b���m��u������˧1��9y�R:�i�O����P�"�E�Ջ��UH��(r��[(D����E<A��JB��̵ָs(X��Z1� �
�V F�2��3�}��Pw��<�QW�Y�;$@Bm�����ݗ���i���&�+��9����P��~�鈢��g�	�5�=��)�i����9��n�����n��~�w~���>��ѣGEv�څW�� �������G�$W���)���@)�g?�7�_����g<O�o`ff��_�]Q/z��.澱x�o>������,���� F�~h� �JO��>�/��|�	f��	
��y�ZH H���x<�P9���=����Gش
y����Q�L:�"�G�J���@���~V
.�8s���� J��plҖ���ݲM7uԚR���,��g�lB.F�2���k!t�уd�U!�����P��I�K��3�o��Q��2/�!�&F�&�E6"/�//wcc�G�l4~�6�sl۶�����3338r� ��q�^���ڵƬ!��v��_0�x�}:%I���y�@�����F����ɫcjj
J�p��mii	۷o����9�<���buu��r�7a��`��C�)ҧ�z$|���� }N3������&\{�ʫj�Ku�%�HP��Hk.UZj�ܪe��*`D�# $t�ܠV�������=96~��y���&RV�\`y�*�C4�9���X#�-c��A�4�G0����E&���3���d��Z 
'wA�e	���A6�6��H���fk�AQ�����o/�
r�u�=�
}p�f-�t���,=2���2����O�+��d��Mʋ����β�3U�G��LJ)��S2xrY#$�������czz�����׿�}��avv_��q�� n��f�y��я~�Z��]�va���Ȳ{���a�i"�����n�2�NY�n�����/��k��_X&��`0�j��bdP8��
�����M�-,�� �ZKk�~�w�>Y��Ç��l(���i#b�8Ӹs̀�4��&���rz�'6�=g���I)�C���h,}�#�w>��}k�7�P<?�-�ĩ}8-.�JE��"�T�X�JG��bߊX�:�͊C[�0Jy�Ø@�(�p��3��PQ�T�����1���ُ��h�X��4?}��z_$�dl!������7��=1:�j�������lWU{y۸P���ԏ��|�N�+^9i�_�v���1b��[����K.��^{-n����u��]w݅��������.|����e�]�+���v��G��7����[k=�p�����*2�:c�j�<�࡙I@*���OX�V���:�rk P�ױ���k��w�y���k$d�Pc��d_W1�qsP^�Hs��9X�z��'�B>*O�3n�W�����r��^�i�/i�1.�̘9�O	;Vi˘��s�X��@�b菚6�	(�I�W�,,rf�w��ݠp��J�W̭ͽ��1�卻��f�=B�t���B����Г�j�|Nj��� �o\��r�n����u����?��y�8�����?333x���G?��ؽ{7���'�s΁1g�q���V�V˻J&I��-�F�� ���~��"Ⱥ�> 3���Gt�=K� ��L����\�e:�n��f��_�/}�K�8G2[��B�,�BLkR
�I��8F���?34��	�Ӓ���U=C��nq�^%H�r��]��B�C��0H`� 75�V#3�|n�\�_��G��U
�1��7�8�F�q��g���_�\Z�7�����4��xIH��J��,�+�I,��UPp��1B|(qb	�������4U�J��{���Bu<��	BY�2C��k��W�УwVVV�k�.|�+_��>�)\r�%طoVWWq��gcyy'�t���'!�2<��υR
x�S��f��믿��r.��,,,�ZgZ��QS����8�=��L���V�amm͛��{�i1��-r���� ����Mk�Ç��O����8�̇��ѣ^s dGځ�P��8��~8}HF*+��V�)���_�~����$]�k�B�!�4�:ĚB@�c���P�8k��q�3�y2�pk:(�!},Җ!}|�-�h�P?�(�
��X5 Sx�(�8�P�����F�:χ���uZ!k-"�<�5s�����ΤTET�~R����w�s��VU���	��Kx�ե55��n�~k8p�ֻ]����,C��G?M������i�#�Μs��W�O��O��sss����u�����Q>%Z���J)�5��^��۔S��X�U��M���h�c �C���Ю�0�.��:�������f�K>��e^H�;�I����T���.�uh�C�[2�q�!�	1ت=��?O��n������3�Z����A!�B�8j"�ۥ�l 7c;�#���GY��:�|~��M[n��*��ۊ��
1VkK�H�>���h�Ӣ��x�[��(��g�V�84zF�6~m��B-�:��ĸ:H�7İ%�M�*�j����4��矏���%8餓<R'�JE8r�Hi��P���".��B\r�%x������#�st: �>ĸ�:(��7ԏ�͐'O�e���رc����i#�R�հ���(���ZV��N��C��Mo��wߍ]�vyO2	p�94�|�`H0LJ!�>I+�AU³j��<�=�kM�줶�$���g����Cs��EO�|p�-� v�?^�8��!u_Ӗ1})���Б��)���JAJ����o3@����NkS/D�Đ_UD���euh���w�
3F�N��Db�ö�
��6M�n��$�������`�m!�K���w�܉o~���K���~�v��j4 ����NU�I�_������V���8+++���W��=���~�3�'���;'��ǖ�,$p���p��Q\{��v�X9��[n���8��.�u�mX��`m���V�4���S���~���1�x��=��C�t�]��>t���q��/�'��!k*K�7�Yn��$�H����9(뼙re[���q7�M�Vk@��K?�R1�N`���]��T���
7��Q�U��X�-c����WM�$�??�{LF%��D�v�.ȥtU
JU�wH8l��&�@�Gi��VM�q�?��˺���d��&=+��x�)�5q��'���~6�8�(���*�\�1:�j���~#�~�w��[n���?�p~~?���o��o��c��>�B��c�I�����7�G�Gؿ?>�����K/�m�݆���}��?�s�q��|�#x�k_���\u�Ux��_������g>����%�l�����^{-v��	k�����zW�eh�CWޗ���P���o(����Ƚ�~�|�i5��+�U%yEQ䵹f��	O��o��/���*m]3� �rӅ�+�)���j� G��X��dܢ+}���}����F7�����m����nq(E�$��R1⨎�.C�G���宖ǈ X�|�C�C�ܽ�D�r�s�/4^���ï�S�먬�>�0��{R���*�#F2+P���q�F��tV(�3����l��?�>�,\u�U�XYF������q�)��g�ރn��}����뾇��Yl߾?���%5����G�瘛�+�p����-<��D�����
 xM��o����w ��juu'�t~�W~۷oǮ����_J�L/�����4Mqx=ö������n͡����S��V
�6��,½K]�q�ބE������G~Z�惵�J3f����
�`��^�0�}n�(�5T1�D'|� -D���=#D#��t�k�h�?C�Ǳ_� �t>��=�����b�Z�i�{IAo��4M)�ug@���R���$�0�Ϡ�ށ(�ak5d� �p�@Y#/hX!�r��86�#(��ш�@fsdy���[�� P1����P�bl��)�&�I�oDH�������<�NY��w�lZ���g�P���:�r�WF�&ib�TF�eP�}l�Ne�P 0$|`�I�_��b�.���CS��_���x�ܪz��/�<���������[n��]v���'����c�������+�D��x�_���������җ��^z)v��|�;�j�p��;��i�Ǟ�l�����&����$薖��Ї>{��0p���O~2 ��O�kV�y�s�P���/����8�S�=�Z�z�\r	�Ї���#��lll�^�mr!�P�ǍI��;��V!�4��!�+���*B����n|�Qÿ́4F�����})Y4����uP��n ��E�I�+I���c���黏��Ѻ�%)3�GU���Qa�P
@�H'H3��u�EV���,w6��@b��w�8d������QJ9�L6�p"�g�s�Z��b���,���P��P���{U����jӽ*�z����.���𲗽�v�B�XXX���<����X^^��ݻ��'?zЃ��¯�گ!Jj��G����i󔟸fx��܉,�!�j���@©��azz�m
kOc}ui��^�;Ğ��y�f����%t:ԓG/�����=��s�����o�o��sp���l��n����6RK=����M�9�1M>>U���Fj�#�h�kv=�x��9�OH���M����\�EĿ�v����Ȳ�$q@�N�3:��#������Jǀ� ��p�� 2�Aiڌ�뾤-�����:4�X*d�τ�}��E@n�1�%S�*� XU��%��a�[>.P.��6�wC�?�%{�����P�fRI�:�CJ�\-F�T�O�+G-Y���k�v�}�s���E�?�|��}�y��Q�W��PJaii	�{��[�����l���d�!S_��Z�4��[��Ea��ݮG��0�$qG:����@��B��ǡC�p�)��7~�7�w�^<xП��� ��d�G��{��V1g9V!����6V��eWՃ?[5wx=d[e��kR�p!����
^�d�Cڡ����d���g-�ѵ%���K0}k;4��"��)�u&�<@�=x�U0>r�qɈLY
VG ��2`���9�1������Q���t�(�&���v$"�2��|(�lhBW�{�B��l�_��Ԟ�����DIs�),-ϱx�h�؝]E��{ �f�Ԍ3�h�����:>�ۅ�nLn:�L_2|�'�0�s���`0���2�ͦؖ��������u��]��/�ܠ^��ޙA�׃��FY�Z��9�'��~���x򏤗�2Fy]��8���C�^��O)��"Pqf7n�Y�Y��%�ῳ�iC!9������te�.�*N1��IRa��#��Fn���I��t�3B,�(b��
6��W>1����Yw��O?�G��;� 9p�Z��¢���6s��7O�]_���~E�j���u�8��^��[�b�!�V�$���,c#��($���䴱��#JfY�#P�لƊ���R~�Z�m�t����#yy���<Q��,˼ǆ1Ư���`}}݇D&�Ou�so��&��|���7��MLOO�2�n����4������o�W�߸1��`�)Dk��0��*o�����>@x�9�����\��u$��~�������������ܦ�
�v�P:TkRX��&t�*�)R#���44ҁ��
:*���/:���w"�������"���Q�f:X�8M��/ј�
�yI"�yJ&B2���\j0Tvh��ʶ/�\����[�z���3C����`uuՇ4��4==��,S�Ą�<B̟&�ɽv(_i��c����7_ѡ&��v��t�QKblll���V�5�mc���ic0`eu	g=�!�_ox=N:�$䅉+I����E�1c�;)�%V��XU����?S���1K����R,$݇���w�����hǧa`��3�CY�� 79r�G$Ϣ�_)�R�:�1����]=]����*m�����c¦p7���:K��Hj`8�Z+X��m�<���ܙ�0,/�sX�")P!]�*����L�Y�O"�������j��x�H�.ϗ��R�T����w�������I5�>4�,MS���jyuc�7�,--�k]t�]DQ���S�5�#�l����k��������%�o��������B���'c�i�V� ��O����|&�����_�m����������h�����i<��K�M2��^��h!z��V�!Ĵ��T�Z4���HC�	v�i�9�}�v.�I4,S8k��X�1��Z��)�7�NH�r,Җn�Rjx����I���MŐgd��,M8��Y`U�Qhd�T�7�i]lo�
�zm8!`0�w���	#41h�C�ę7�P���̈��C��p��O �;����(�������ʒ��Au���ן���+�A���o�)��ӻq{�(�|b���H)�=w�h��LDy��w�k��.����������>zfE~3U�����;P��X؎���� '��F���l��G-NЙ��lg�^+K˾�d�"��͑$��^4>$(9=R��?;����C�<~>�-�%?h�ƚ
�9�(_n
��Tw�b��7�rړZ�;z�� 3�d� '	��2k��8��Z�̓D#��Z���d�5`�;S770�@���%�i���Ok!���3�P��{,Җz�3dQyO�,�1��0�LR�/�+��T��fPp�����4E�~��g�0@��{�:��d�~�H�@�2_��d�DM"0B1�����˪z�7?ȉI�k�����n���T�z�ݮ���}�<{h���Ԕ?�jcc����`��ѹ�T�^�~����c��(I4�M:t�~��qꩧ�iO{�_#����������[�c:t��˿��~�����Ǔ��d|�ӟF�ex򓟌/��Ȳ�zԣ��o~ �G=
?��Opd�(��݋N��i��9@ߜ�GPfޒfH�#��ʫhaҬ�"�4}��3p	08p�vqj�'���� 8�������K
�td�8Fo�?	0�.^d�ǑU�8���P����2A�`�f�c���{��w�'�s�TEŉW���oSӬ��.�ɋ��Ҁq'a�br�1�� ��o���/�>�2s��CDJ�R��v�R=eUy���T]��Bm	�������64���G2���GH{�������§8� �[����=�M!d�'���m�p��Xk������%,--aaa p��QLMM�Z��L���oll�?�fgg}��$I��}_�����?_��Wp�w�S�O|�8�3���?���?�����s�����
W��x�������/�������/����s�N�/�4���i�'�����/rT-\����΀)I2��e�� �D�\�$D���#>�FA��+Vi�b/ѐf�v�!�9Ӏ6�#�#@iǒ�J�&E�HG,�(v���жK����|������z�U�Oa������s�� ��xɌP�����;.�"�B=�a��`C�d~C�7z��'��9I�!�V2�P
1~z�&/���"��!�_5���+������n;v��g>�\y啸���<��;�����l6155�{�����R!WJc:�����}'�p��o۷o������i�m۶acc�F�#)�/c�Ν�袋��z����t:x򓟌?��8�����?ߟ}��>����<>|���x�s� 8������똚�B�x�c�N����Y����|�����o�T%�%��1�c<�sHC��_��*����t"��{$ؑ�q���͕�p����r�A��;�J3�;+�(�(�0 sUT�_����ܮ-�u!2�*�JQh�e�2��[� �(A�;�o���n���8 ���A�b@7 ��k�1��"Ms���s:����B�܅R~��J��'0R����&��[���!��PGF.0�B�U!EY�P;(��k+˘j5Q�#��h��u4j	�I��h���ԓ������~��೟�,��:�mۆ<�1==���9�x㍸袋p뭷���+_�J|���G������6��Mo�`0���l����K���>�1|�����*���p���ٳO|��n�qꩧ���FEx�c��=�q8p� n���=��o���� ~�7�|�3q������>�����+-:S���N�'׆Bvm>Un�R��b���S��f�Rj�Tց���LC���0�_��JBD[X-qß��Y�0�F�)d�En �+�J���E^�ߛdlﯯ]��a������|����8���K���;I�фzIPL�H�:�f��vy�C�B�Zf6Bk��^�FU_�3���:vRgK��U�a36�& ��ׁ�7]�����I��ǟ��%
����ƺȗ'�|2^���c�޽��O���y=z���9EnQ��O��^�:��s�W�)����<��;���;wb۶m��_�u�ٳ�~�|�#j��0;;����{���U���=�� SSSX^^���2 x-pqy��n���ݻ�Z,--�Z��k���ߏ�|�#�t:>��'��f���P�Ch8�����帍�r�$��g�ZY�|'�q���=�X���&!�|VGt�����w]4T����ȓa�E(2�)�xhF���&���1�A&���>��;[��cw�]�+(��-�������1mKQ*-�"@���W�e6�@T�Q'��b��!6m]L�a��vp����Q���GR��-��!���r����e��$=�$	-r��H�9�R��g�~���M7݄}�����o�i������cvv����x�{����k�z�8묳��o��+OA���G?�Qlll�����Z����9���������׼y���ѣx�s��N�����
W]u�G`ffƷ���bvv�Zg�uZ�����F����(B��zƖ�u<����mx��|9��Hb��L�d}��<�8�a��O.{���^���;@��dc�iH0M���C4R������@�rU�C�����+%ϟ�)YgY�Ѿ�RS�;'D)6@נ�[wJ��hh�V�F�^���4E��?�&�-c�O��Ǭ��sp▃1�3��r����
�<w�~I�:G�$��T�rFk��)'Kڕ.��>%i����y���5�3p"ƒ�AE���H���U�C
9:_��.@�������>Z��_9z�(��.�n��Vl߾�·��-�q�Y8���q�M7���{"G�L6�n���}�s��׾���㘚���Ç���,�p��\~��سg���p�^H{
�4E���`�B2:t���'���	'����ݮ�}�o��o�ַ��Az.�����$�/}�Ǭ���9��Z�D�!f̙,�*<N��4.�8���9:�f.j��M��P���)���6��I
`�2r��g��Hj	L�1H3D&��'/tm���]��� �P��~r�=i�r�:��:+�5��PVA�}�t� ��k�@cD�s�sF��B<�M��
� G��VH)��GH�F� ]hmя��PG]t��X�T�&2���K�T'�oNdҮO����249��9(Ǥ�*w�����L��<�$�1��$ O���'61ސj�c��4y. ���4�S8�����.~��=g�q��6�����t������)$I�7��r�j5t:|���5���7sQݒ$)-�+�<���_��xzzڻr��m��o�6��w-�IHn�i�BG@nRd� �F��T{N؍��)@�&lR��t�h�����6<����"Z���B�֎R�<�R�	r.Ɨ���"����6}s�C�?��cH&������d�w8�s�L���<�tJB�J�)/c0Ơ97a�ؙ|��R7�u��8i����:������2� �7�Q��8��V�a����̙�rXgi�
J�z�Q&׈b��Xh8>uW_���;5d
q�>�u_�Pr�EយA{�뉐�ÿ�]NX)�IG�Ù+F�A�T:�B�:g���R�� ']U?���LR�HM�Jˑ���f��[n��x�;��<g�}������۷o��Ν;}�v����t:%�C~�<n	�n��Z��N8g�}6:����8t����gannG��Rʟ�����n���2������*���-�IOz�7-eY�l*�����3�<_|1�r'�8p���K�h�H�)�Ǎah����d��N���$��8��B�JC����̸�m�ό !�h�ȝ�5�g@Jn�&/��l�"����U֠�d��_>J[�d��iJ@ 5s�`"<I��ֽ�ζ�<J�R0��t&Mjz���.�$���B���
1sJ�� ��a���W�C>'�������׿��xғ����et�]�y�"V���4C�OzC�#�L��?G �*�o����ָ��q���cyyY�y�{��^����-�<���S�5�����,VWW}4��/��~����g~~�#���i�z뭸��K�o| �}R�%�&�}+w�3DkU�h|\C4E�G}��;ӥ(����:�1��V�_k��c�U�b/�!��a�p��z	��&��P��.N�^$n.��v�6�����o�w�'QR�l�A��E�q��̋ۓ)�0hq��x�!�m���,���9a��2�=�`
]�4)B�*�<.��d�]ޛ$4B���~���?���v��qnllx���7�w��~"aLcA��!yܬ��z���� ���ؽ{�۶m�E]���9��1>8Z�V�`0(1k�1��'<�o�"��(�077���)��u<���Ν;1��Tgڀ�ib� ��5>n\��b�!�
�k�P!�JȓF.���rBz�̓����$��c���iAc1���Yf`��WhdJ
2�Ja:����a��M�9�]�C��QA�<�bG��o���	����i�;a�>�	"v���pC���>�O��a��P�!m"��8��Ҥ�*�%�t��,S�m��G������h4�����%Y���h�pdS���~0x[0!��`�>�Q�s�3�@����W_�������D<��OƝwމ`�Νh�Z���&���t�+�_�B ���"������l�~���|Y���8���7"I/��A1.<��#��f/���V)��������ϯI&�x�<��e���*�9�"X��b@%�Ո�.8ڐ^M>'�]H[��w�?qKY�sJ�G0}�a���P� V��2m�y�M��)������#ymf`%ӕ��$D�J[���'��`<�OF�$s�8�%����.��ғa�;|�d��2�N�/�&gdy�b�8w����S�}�ӓ����E�S�6}򺡠k�Cׇ���*���p�-�x��������?�y��mt:oΡ<Ik��AD#��v��������~�u�]��'>��������133���n��0��A�)thmE��8dXE|NȹB��@%,QΏ*Ms-r�wt93��h��kR�	%z�<�H�� y<X!|�_5>����V�ͱH[����R'�F ,L� �����яA��X��V�0��lq�"��� ���p\r��	�3[�`�`n��1	m��G_�L�=1MWw�QK����8�??Ę��O����������4�4����7�$I��x��Z��j�]���Ez�����*�8���mo���<VWW�׼���OɬC��E\l���i��e/C�رc~�����ضm��֜�H�hKa��<���Ic�}�m�60Nr\��])�7�Ə����C˜>�4q��[U�|H+�����/����R�9����RƇu�y��u!e��������t�����3��+��$�!ڷ�-N��p|0�ø;P�z��p���n���"g@�0,�
*��#��a��a��B�C�4�Yfkg� 4Ah��t@�u�3w��$���&"t�I���&Hy��Q����|��ø{!T���6�͔b �I�A}L'`q���Z@������~N��ɻ��C:��LF�t�=�w��t�]���t:ؿ�;e}����f*��~2KMMM�]�J)<�)OA�$X\\�#�H�ر���X__w�bb��k�Z��]���5eL���4B�U�9���@�o��R{8�ыt���BZ�94�7������ϒ�E��F#�r�6/xC�(c4���,:�+hD����Xa����H[��v�:���~�A�yi�2Ɠ.g.�b�m��%�8�u~��F
"]G-i!�z�>��N첀�$*�;��3\"RщH��zi����V�d^�����@X�1�e�|� ��A}%C�r�>�B�aYg�*�˫P�� ���\��������q�4�F����2��i����CVh��ݮ�l���P�t:����>��NQ��`Ą�puڌE�{��TZ+ �@}����C��>���{K�{>�|ܨ�=��B4C!��d��6@�s����tF�cK�)�;��8�yF���].�9���R>��:�'>h��y��=����������L�N�`���)���+ޯ4�d��H�<M$����i&�"$���ɟ�������bӗ̎30����@�Uj*�G�I�h$� @��85*�r9�ɼ�f�?��O�u^_�R�Z����Ky]��P?IMf���M6�v�k�?]�^��	G��i�Z^�ѽ��˿�'?�I�!��	 �TH�������7ވk��I���{��7� �n��8p ���8r���ߏN��! ���<) Ǚ��Ԅ�gj��J;71-�r9��eK�^�^�]���*�k�!fΟ��$�!f�OG#M��!��̒|��;|3�%��B��ͅLa��u�c!:�?��ıJ[���.�E(�b��EB6�gP�؆��~����:�����OV��Wȉ+'W�P>�B"&��dUnl�$���!�r��H,$�I(��I[�䳄�fggQ��155���illl�S��⹵.�!�v�����|�����W��O��������ƽ�ދ+������e�����+��u�]�׾������q�����x�ߌ����^c 4Z�		=>>�e�����U�D��?ћ*���4���-�V1S	Xd�9@B�j݈�6��;!��xO�QS�<�!�S8?{��`,���z���2/+���."{���ϱH[��K�b�z�7f�8���z��wr��3N���9�q;�=s^2}iR��Ѥ��L�Hf �)��>�*��߫b���q�B���u��F��,�p��7cffJ)8p��¥�V4�j��?$���ammxի^c�Ʃ��_y�LOO�V�a�޽x�ӟ���y\p�^x�C�V����9<�я�޽{1��?w�}7��w%�O��Nm14�g�/�`�t�����B��y�ߕ�R�l���m�ϟ	�9�����ȅC�G�>ֺ������� Sb���Ͳ��P��~��R�G?
��P��<s�[�	��L�����ίu>��9�1�ݞ\t����F��u+ �b������s�b�"��1�*$˙{��b��2���5��<x��84ȟ��ܱLRpR�t:�����w�;v���^~��8z�(^��W�1�y^�җz~k� Zk��}�C��x�+_	k->����i���i���?����><�ĳ��,Xkq�=���~��E�����<���/��"c������E�N���華#F��9������� O�.KL. x���;!�����h��Hx�����Zg���\'	Q�B&Qه�ق/�k�%��U>�/��In�ZV+�y�4w�:*�5�`3���`~��N�Ɂ��P����_aX9[~A�QiL�o�r�B��=��X/�n�J)�U��T� PS�(��'�jB�R���%��BRiK�`��G��ݪ��T��x$���'����Zg�������(LOO{�|�1�s�=�������q�=�`}}333���wމ~��Çc۶mضm�wu�Eۯ�똙��c�X,//��ص�5wVr��}�	��j59r�u�v�N$������d������K�U��w%��_e���s��P�Bc�K�/���C�E���S��:=���Q,C펵�מU�>�Z�0��$v�5(��7���sGn�?@�=��?˴���h�R��3�3 ���	e�N(GӀjwr�2�8�!�J�_��h"�;!�!'���8^=+�F����m*���ǤIz��[��|\ۭu��ܹ�x�+���aff�^z)���p��7czz�o�����f/��Ev�څ�^�{7�#G���N���ٟ���`ee�3u
�@�C4���2���P��0===r|���P��P���=��=άCT)%ʒ�Ù�\<�c��m�-�����gd�BS���+D�����R#�m�xO+(�]��f�s�����,i@C'����4�醛fT�)̾Ú��4�����i�r�6�T<C5�-ɞ��C�% .�T}�k�'˕�CDM���q�vHf�G��B�}���w�qH�\%�BeN��B�B-,//�ȑ#X^^�.�qczz�^{-~���\s���}�ri��W��w������tP��P����O~�y�kp�]w��x�j�$��,w��=m�"�P�R����� �H5d���U�Q2q.���+=H�=���pwIb(!M�B��^�nx���r�u�m
ѹ\���/�/���/���Y�'D������d[>���G��� |~�x�Rã!��E�2��h��s �����wy�_:PؤF[w�I�L7F)�Z!6� O#GO�0*C�&��a������ ۀ�)t��Fd��<�C�&�(F>��N"���,�@G9�	�$�&ǈ�������1n΃�~�_.JqT�Q����o(��~"�J�0��'�*�R�x�|�ѽZ�z�3�Z��~����w�q8��s1??�f��v����5 ��).N�� �<ϱ��cLi-�\�hAV)�<��y��C��P��#�i'�p~�q��1�Bt��T�Ӎ��|����) Z�� �c��P�c���?7�P]�m�2(�i�f!�q�O�HȒi��H�7�JZ�������x����!�}Qm ���Y����$���"D��D�jX���<��][q�!�}B�ZX�����l�p�6��@[h�"D
�uh����i K��w���3�l�w�����H}fu!̤D<B�b�l�MP�	��	3�2�8�&�^�D�5��R������O�*t/�-�#Ss�ώs�D���|�����&�^�;�~�4�����8�3��7�i��k������h�Z��jx���s�9'�x"666���9�y��ԧ�����;�R��%�N����yAC��a��̠�����5b��O܅�B7��Q=P���d~Ĝ���8�GٷUZ���]q[�縼$�B?�e���*�#�L��s�ý���Q��-6��)H�B)�b���cû�}���I��Vx}��z=�U��e����׬�P���1��E���~�e"10&�1É��)�����yQ�m��x�:!,R�H���J�Xe"
1H)(y�r��I5�	��6P�q�CχTQ�����,)�B��Z-�z=?1��/����	��h��k�������k_�:���+�5����[n���^�������SSS�C.(�%b�I��yP 8����0P�Ւָ)O��)�Ɖ?#ˑ^-W�Ks����gǥ�z�̕U�P��r����HU{�Ϻ���*(�C��a1�p)�>�x?�o�6�-���p�0�%�*m���z(� D�7����T(f�@a2F1�k֖���?�QA1�=��Z%PJ�S&�������'1�P��PUm�EN���q�C���ph��\�{�Q�S�fggq�b�޽%gcVVV|��F��v��z��{�sss������v�h6��dD{
�y�۝���|,�5��%��kT���ȹ
D��K��f9P�i���ʕ�;���gCm�s���y>t�.ER1��~�b!��O��sg�6��
E&Kk7w�,|<~�K���6�.'-�ߗ�����e&�,���]�׾���b���sJʸ��BG@6Ȃ��$��a�#m��Xes8a%��֩�#��f�x!Q^xuM�O�wx����\̈́��B�D
�
�C��d�M���b<Zk'�2<��υ1�����C�����x���0==��z_���Xk�{�n\t�Eh6�8t�>�ݻw�����ajj���[�VVV����=�����Ck�c�P�OK�O4#=|�6��)�"�t��O$�!Z��-ˑ�+��`M��1�A
�*-R
7Ik� y��C��Kk�k$ƝY)w�a%��E���Z!��͚���2�����qYS�Ԁ��;�v���]<nr�q��G���O�2󎋟R>��1�p��#<4�@�r��JH�BM�eJ5��������	���=��&��E�	4�!o��~�I���v�k��8A�� ��"�\�$	�=�W������>���%\r�%��?��۷�����z/���5���`ffW^y%���7�������?�����ȲW^y%>����n�;��|�_D�V�g>���}���!*�]�׀������f?ޟ����h��8m�c>r����A�}�B�A�����U�5	�5��ҫ��{J����?�/Bt��u*��ZP%D"�s,���/��E���X���3׽}N�NG� y(��'�{ǚb!�*����f06l���`]"�����<48���(���BJ!�S��8"�ͤ��U(+�'��/�?If.y�����/x򐇠V��iO{N<�D,//{�K��Y�d�!��N����I�`eekkk���8z���箻��O~����'yQDP�6��������hD2y��������#���bH�����ҩD�!!$�����/�T��n���*�G0���n<k�����Tsg�K��N���h���cpm˘����~s��=�&�L%)��J)h�KZ��(�L!�/тD�I��[&���������#�e��ه�OJ�I;.�ty�g��,��7�Zh�Dh�����nccc�FQaqq�������]���%/y	�1X__����(��������<�fO��=�}�K^����K.��%/y	��>���|���_�����!s#%���Lj�d�4��4�KU�!4&!����G�y�d� ���:�hJ�VY�9�{�7�0����T��/���C�_h��١����Z��*0!`��*-����2�f��F���(V���f(P �P�3i(���"S���"*��+�`ld)r�AY�$���M�] D��h*��6W^�
�f4`d/䈇�%�k�hB2NN���P�n}�EQ J!s�j�,K��Є�}��MB�����A���T'rc�z��O��OMMayy����z��µ�5�g��(�1>?B�T��o4~Qvjj
J9��;wB)���l۶�ӂR�o���N���������4��Gd�3�F��9#�s�����ƚ�P��q�c-���=__��С��rz���{*�ʭ��#m.�lH ���m�����]R�eY��º�Z���:�!�-42(
��]�6�0HsD��	�i���9";^F��Z�8A�����%��*�E�[hӀk[ZY�Q�Zb26���T?�܁HL�_�:�#p��b��g�͓ҸwB���еII�Ҕ���rMD�[��g$����}N�����gH�
KG���annQ�^�cff�N���1����,(�(rg�Z����:/�v]� X]]���Z�c�SX����e���?==]21��)�՘p�ͯ�q���'�J�!>?ǕJ!mP�_�6�q�m�t#=���W`t��Q��zO��Ɔ�o�� ��X��}��;����ϛ��{ �Q�3[2��Nt���g�[�VJO�����C�����al�g���<�V9�q�e�B�;��i��h�@L��׽jҎ#b9����H*#T�S F�3��'5��)Im�TU.��<���VWWq����Ùg��/|��o��amm���w�ԧ>�������������W��;���k��F�c�ъ��w]����A2Z�!��e�����v�n_Z����� WVV0;;k-666�}�v��}�xuuտR���s\U�P���<I ß7��oeݥ�'$��9ǯW}�������� �Ykh�q��`��]�dXc�1.|��
�V	����*�5Jq���ܱ���Z���g3 p�iː�S���-�S	�UHt��ƥ��F��!F͟��R�,�
��eUM���R�e�6{=�P(��Q�,[2�>GW�6I����g?C��������jt�]�߿���wq��A|�{��7� c���z|�3��jB��Zt:�Ə���3z ޼��Vtx����k�G�G������}�s��˰���o~���?�#�x��ַ��K/���v����8��3r^�=�B�BΉ���&!U>?6�Bυ5�ːW��k(O���U����g xs7�8�Ҷ6�u���i�Z�nH���6��<�� ���M��0I�H��P�b�t2k�"@Ù�������PPȡm��1���l�Vƅ�d��>�,QJ�#QO��l
	ѐ �>�u�b�!-�כ��w-[;?\�#��C'_�}�ݸ����7��f�W�W�����'��s�=۷o�I'��nםM��g<���1??��(�^�{�H�99r�WJy��ҡ���;wBk�myy�3�PL�<�}���k����8���PJ�8?�fb|����0�>I||CK�?龬�S�w�9N�U�dY�βOB���K)�Lй�`��
��K.���������\3}B��d��p��
0eWw��p�X��1}'����$��Z�H���G�<U~��|����q5!��!j�����yޛ��g�bhrLb���0`tɅ=ɸBu�kd���׾�����x��އG=�Q8r�Z�����j�p�q�auu{��AE8x� ����s���W^�/��x�3��G?��^{ ���DH�#��orפ�ԭ���׿��?�{���G=
Zk�|��x���O<+++x�k^�?�����ǹ瞋�{��;�@��~����}B�x�����UU��,���GH8�{!�#˓�'y����>����:��뭉�^Y��tY��2�l��-3~X�}��I[��KcVbvV�U�
f02���|c�П_�n ���2�����L^����@���ǟ�>��ke;1J�U�-��d�!�M	���:�we���k�D^�!U	m������^������ѣX[[�q�����=z�f���8r��4Ł���J��r��*�I�^�����R�ķN���o�_|1���333ؾ};��::�������_��_�+����2�;�8<�����*��w�����$�b�=�� dݫ����S������7�yK�g�!"\[W^�b����w*��"X��Le���yWe������-׿�U��CTx=G	w|#���*�|G��A�$p|�W#��D�oi�Ǭ��#?�l&'g���iï��u�j1����		Y;��Se?����&�=�Z��3�8�5�1�R~�����z�غ��\x�8�Ӱk�.<x�z�fӛxF��r�q�#�P?�-���^�����عs'�����SNA�����h�d���g���(`��n�ZX[[��ݻ���d��x]x;d�c�6s&/�x ��4e�T�i�D���B��*w�q�I-��FHpc`l ʧ�����7��w��m����Vѐ_��A>� n6m�w�f�Ql��&tb��dj*1���-VƑC%�VƘ����D0ykb�T6��)h4a#���`�#�s�A��,�ш�4��߹ks�XG�P��H��q7bDQ:�Nő>�\B�Ee"8�|�:��7h������*E2�*�Du�������	%
E���[�O��������W�
����177�~���(�~�����ݧ���|�]v���z������MRC�gjq��ߖmܹ��)rk�~��Q&�c��X�߆^���i4���@�ex�c��?��>����2fgg�7��zիP��q�]w���Z����S��?T�|�`v)�H�pZ��A`�wF
�m�ᐫ���CGsg�����Q{9�Jp��]��|A�Ӵl[?[� ߀A�QD��K�'�u��ju�V�� v
:n������҈�u�lJ�0�#��A
9"��`2UC�5�����@��c��Ĉ�ȁa����+Hkhk�Z��c�����u�����&�cHJ��!�T�ډH�&,B!ՏO��rƩ�!�$�̤�Q6_嗓��I�q&�Y�B>�lB�����8�g�}6�����>�1h6������Z�����h4�$�����t�n��w�^�Xk�����>�_��Z�)�3�P������y�y睸�K����Ϙ���{cc�N���u��W\�MT
"�cl߾?�я��������{�Z-��m�H��L�#�&�ƅ{�`����(�_�3!TZ�M����5)I-Sj�$�x��69��}�Y�ڒu�����v�ul/�.1�J@M�.W�*m���5�~s�Q5���a�� ��uϿ z�_)w V�"(�â0)Y���L���( ���-�H� s����saS���PUd>�=��чƄ�qܤ���*Oy���`qq�w�Ƴ��l|��_E���Ν;���~��vVVVp��w��SO��wߍf��N87�t�(���D��/��7Q���6s�n�-��Y�c(�;��WW�1�9��O>�'��N:	�����$I���s��\�D��}R8�={����h����M���%SP�����'��1��ǆޕ���M�f��I:�V�?��N&�K@�?��g�Ot��},�۰�5�M�B�d���3}����s>��y�/��p��f�fӖ.��q��h��A�J&�
)
k=ӯB�rPY!&ˉ�� 9QBd��N��|^�3T�H_T$�\8�ZG�|,Bm��k��
	*�(�BǸ���7�W]u����կ~5~���_�*���7�[����O��{������}�Cx��ߎ��U�رi�bee�� �fӗɵ��EU��������i�bqq�/6oll`ffJ)��v���WVV����>��x�ӟ���;SSS~7��.�3��I�?ef4J���G.@��-RRW/Y�*M*d�D�L����©
�h>�=�}�4�҂�����jc������[�ђ�
N]��hGB��*m�5��4��>�"[�XDS���b���u0�<���A_�,*uS��Bj��U�O��8!�/��UE�R�˶Q���{��;�8������ۇz��׼�58�S�(�s����t�'=	������{�E�$>����>�ԧ����I�MOO㦛n�'?�I<�	O�/�z���ݿc�,//������<�q��Hggg155�o�ozӛp����U�z�� ��˥�qRHs�"���^����7�U)ԟ!:�
�l��9���$���:��V��Xc]4 k-r���� �f�Mz-$T���	�<e��>�;�*m�wv��G�y|�II��~Ռ�����2��膜�$J�yK���'�VnK�w7�\8Hm�������������.�͵�$I���>�G�<��3����;v������2���gAk��W�W����Ç�3���&�&�"����̙ ��U��'Ya�9z�(��ك7�������Ç8o#��k����^�� �N�/�6���cffO{���=���X__/�n������*�1B�<0\Ն\)C����hs� G{��L���W��5����������VP� f�P΁��o�fe�,؜�v�v8����Y�k+u��L�׋5�B4|��ȼ�p펏���(�jE�A+������m���6!F"�*��W��<�^!��BC��4�ʖi�Hm3��R�*c\��(�| ���uh�Σ�����H��Z%/r��p�U���@��W���l����bjj�3♙w�qH��z׻p��A\|�Ÿ��[�}�|�#������8p� �4-��Y__�'~�{�ؿ?������ت��^x�b�Kڗ}��?�~V�)��>d���8��S)Gb�
����yy��/��]o*�<�
�{��ӫ����	�jX�+j�}>�����TXk����@��>v�z�7gф��\A�,���#63J�Z���oȇ���qD$��l"4^&o+�O�A��I�1)�x ���'�����I��+ԟ�b�U�?K�Og���+=3���:55���5M�l����%7Z�~��1��3ڜE�x��.�=���E�}��ރ�k��]w݅��U,..���f�	�5�9�N��5>�����/����ݮ�k@m�%�/���X�o��U�G�y,�����U�T��9�=�xU�5$HB����!�"=jB�%�f�^�?R/��|��X�-��E�`���S�����z��8Ϟ�I(�űF������ZJ�8���]��)[cǔWέv��&�R�'�,5E,r�р$:�0���YRŖL��C̘/hӵ* �>' B���+�O_�� &�= h"��*9a� �k<q$���3*>q�s�Vk�q���f��z���";�1kkkh6�������=T?�<MS�j5�����n�7YkK��P?Q윗����v�سg����̟�����WQ�����Ӟ�4��/�"v���ǲ�j�^���Q��O&+k��f8MJ�G���\r�x<�]� �6y��eNyp�*��u)F=+]���\H����h��<���yһ��=�Z7��b��(��9�>fff�(q�Vk�����Q�i�7�h���sıF���dd�P�r�3YR?����%&	�1F��[�
/vX(k���r�_9�R
�� 9"��(��8����T���$ڸ�C�(�Ǥr9�9d�B�D
.L���D�����Du O:)�U��)6�ۓ�9��&�����kkk~a�1�	����Q9m��MFW��jaii	SSS~0iI�x!������`0�i��潈Z�666�������}<�я�n�����d0i�猒�{i-�1��"nh_ϟ�2�KZ"�<�.��mѧ��k�@`�����[�e0`׆���1�~��	�HM����i[���F����̼�$��X�q���$�!Se"������±�(��(��PN�j�	dX��"�D3U���)E�G���Cu�J%ղH!�S������H�#��3#^�̯V�!�2LMMa}}����,�|���5�z=��	���{��������8���tiawvv���l6�j@����}��}w:��4�!�0Y�h�VsZ�1H6??���u��ul۶͇l���A��ƶm��n�q��A4������G��\�H�����3��
-��h��Z��C�>�o�ي���b�	�P;�KfhIo$�I�:�y!��R��P�$�D��:�(�B�ı�;6U�:CY�Wh�s�E���6})�F���W1(~�3����$X�87yx>!{�I2�P[Bu�z�{�zW!5�_H`H�5���P�1H��:h2��?�#�������g��׿_�җ�����x�K_�뮻W_}5^����{����< �G��K�w����+��7��Z��g?�k^�\w�u���E����u�jvv��z+����������t�0b$��{�����<�4šC��|qcuu7�p�,Í7ވ�z�p�]wa۶m~Q����H��	�L��$i5�^5��Ve=��������#!���7�C(���w\I�.�	2Y��M�2�x��=���x
��9��˱H[��ݠTŔ�/���q.aZ ��a�ڂΓ�-,�l�)L�F��a�Y�c��Ee_� ����������wB��8b�D*���hy�2�ʅ�1�������}r��t:�t:8��q�I'���`nnqc���سg����Mf�v��M9�]�	8p �:��O~�����ކEh4��w��}�C��[0==�,EZĵ�^��/���v>��O�o|#���q�W�-oy����o}+>��Obff���'�׽����;vxaG��.t*��I����k�Vi���*�z��6)�I n0���zθ~�������Zk���\W
�J��la��Q܃�j���>��?.1 q�� (=���JkX�S)��L��W�d3	g��K'T�'���/�MD!a3��!���J�p����W��Z�O̺��p�UW�~�������x���<�q��<��O�9眃,���=�F��v6660;;���9 N�9r�v/~񋽠8����w��Fi��P���Y\x�س�x�w�y^�l��ޅ��l��l�^���O�S��w�q8�S��v1==�]�vᬳ�¶m۰w�^��͕B14�M�×�(��ȋg�x���1=WE�|�$��AB��EN;@9�I��!����yREO��|�~�5�_wU Dߧ��M��]J��<-�S�7B���p@{�Җ1}���;��X혲h䰃�9�^���Ƹ� !�����3���PhZ�:A�����/'�aR�2�c���>	9Q~��/G)狿s�N�q�����+LOO�}(<�Z���;w�o��o��~�}�{q�buu�z_����O|���q�	'����PJ����h�o��o�o|o}�[qꩧbff�z_�җp�W��x��Gayy��^����S���ս��j�3�{�����dh�5S�����#*>��S���'�Fߋ�q$���D3`^Ԙ`�8A0	�<Q��AԠ�t�ݷ��g�{W����ꬽN�}.�7�����{��C�����U�V�3���������m�6���<��v�����cqq/x��q�y��P�^x!�(�E]�(��j��{�n��_�B��/�"fffp�7��O���8���011�sH�)/b
2��d����7W�%}��!M�3F^Y7N@qQY2�2 C�C^C�^	\�� >�" ���)l�e v��G�M�S�Tԟ���5�԰�;���w�7?L�n���3T��eX��텖���� jq�/�Jw�\��I)��$V�.��h�V�$Z(�@�,%�N*���HC��eH~5��9*�V���ѣطo>����SOţ�>�Z��,˰�~�u�Yh4زe �P��r
.��B�C;_i�`˖-طo�?����C������
z��]�����"��yf�|��عs'~���* �믿���x�n��o��ư�����QdY���9taa�F{�����^�w��ݸ袋����ذa�_ĥM\|1����?|p�N�W-����A�x�Z��2�S�6C�Ӥ4�pD�����!~��_����c�E�	P��*1�Z�����
L�% �܋���l[���ؙ~�(/�X�5c��ux]Epq�u
��:�`�� DF������D�����v�H2�0�up/I�} �U�P���L�Zd���� ��1�i�n�p�6��T��PA�>����J������OtAСO���ICCN$9�9�׹�4ݓ��:H��&�QMH��IR{����(��~�z뭨��8��
�"M`yy��m6�8�sp���cnn�^{-6oތN8��͟z�سg������E�:�,�}��PJ������f��s X�1�n
����8�h4x㥗���zwQ��9z�(�ͦ?������%I����cjj
^x!�������?�)J�An��Z�F�
�	o�,��#��7�;w9}��
@�����&h����3Lz�U��yP_��==K�p����UT�Xw��4�J,����IY�8ۼ���@Vk �5`��T
��m��H3��Gw�`d�5�Z��Mk�Q�eDH���b(��5�6T��/�V����������5uٌ�q�!d*�?>y�T}�O��rs�!m�YR�DP�P�V�;O�~���FBL�w��)C]! ���	=[Uvha.��iNr��3��ӹ�9|���Ə�c��H��߿�z׻p�7`���h�Z�4+k-����o�6���Z�FE����o����SSS�ߞ�������x���	SSS>���=z_��p�u�y�3-���?�3n��F9r�f�3���Q��=-V�z=��w�֭صk�?`ii	J)4o�/Cw��e���~�N�r�j�k���V�yo��<�ϯL#�|�3r����t�<�ցH�O⛨
<�	�P_�����;���K�6=�U��:�s�$ÐBG0)c�:G@j�ϋ��]ܼl�P��d~5�1An�����ge�)_S�#SYY����^�'�/�f��_U/���$����p�)��-oy�m��c�7,//㤓N�W\�m۶ᡇ�[k�g׮]��˰q�F?Qz�������lb˖-XYY�����oK��³��l�p�	��S���Q��z�3�N���,///����x������i؆|� 
ͼ���8��n�:\����+��g�q&&&�n�������q4�X�!G�_�9eC�9�:����2���:K� �H	-��^�ͅ���]'�?'���n�SIibQS�X��E\⸎Fc
}�4g��}�m �B���
��]�� Ź�E@�4N
��KH�yt[Q����v�+�d�sQ�.�+����/���,B�LZs��24,�EN�IW%h$ї�_5�����3���F����/�o��o�׼�6m���Z���z��v�>�l�ܹ�#*2#,--�QJ),,,`ll۶m�AܔR���D��h��Ů]��<;w���Z뵌��I��/��8�����[��Z��$I�o}�w����
:��+S��Ui��صk^�������è��n�4���.C�|\C�a�{&�?�_U�d�U��on�a'x�!�]VGَ�:r��A'Ͽ����C/�p}} �n]2h���@�ꛆe�UZ��Y�����'F12w"U��X�0�Gݜ��@Ҥ��y<J&?5+ߝ�R���]8��F��e��U��!A'H�W�L��2f[�,�ow(���i���2"���qlڴ	�ׯG�������.6n܈��E|�k_���ߏ��q�z=,..���b||��?�a�˿��(����e���J|�C��⢏MO.�������[��׿�^{-���g��������;������=���Ǳ7��_�;v��5�\�w�󝘝�ſ���o}+��>�t�M����m��?�3>����������/|�^z)�8ƛ��&�w�y>� 4b��!����\����O��˵�a`��#�h�Z�/�1}�马�P���A��=U}��F ��J�GMX!M҄��I�&�[AcGⵞ��ǚ���������AD��&�N_�r��!C��h��/��W�{'3���\�"a�'g�T^C�������"F����'�TqC9T7��L c��m@qLɯ~Ϟ=����}=z��s�?��;��	'��?��?�1�>��7�Xk�����{����?v�܉$I|x���?� �5�Z��F��^��MJ���o�>o���z��͛q��a<��O��ݻ�h4���d˝�����N<�Do6"z���XYY�R
��-[`��}�݇x G����7R�����
�,���>1
�Uf�yH0W��j�����.��4,�)n��@��B{1�v���Ϸ��24�ҰjP�p�]���9U��E!m� �Ҕ~Ҵ�L�v�ȃ�5j�f�4��C�;AFz�O�w��w��Zeyd�\%d�Z[�J�;bp�E�L_y��y��*��M�2�N�C�e�JM-+�ߗ�)Ԇл��R��̃����Ӹ��{q饗����e�]�������>�1\v�ex�s����m<�2�Z-�p������������t:ػw/��O�?��p��Ϊm��رc�8�=z���g033�3�<���7p��Q�{�x��ߎ��Et:�>��h6��t:��_�E������C��B��?�a4�M�ٳ�/���e/�K^��_�~ �'P�9�?ԏ�F�X<{pH����LC6�e�Z�ə�cHg
���C��,3(,3� !~2�j]����{"iCk����#�Y�+�4t-�6�aY���re�����a"��[�R��a�걦53�P����ŏ �F��#}�
��=1��3^C;��oyjT��%�p��v^�H	\�C���"P��B�r�+���*?�	��Ų�~Ȍ0,)�<ä���{.N:�$c�u�V�������O;bi�*�Z...�;���7����G���;��<�s���f���8z�(fgg�7�7��'?�V��/~���?���9�z=,//��\j3E�$7�4M111���Qt:��̠�jA)��۷c˖-X\\���4�n�����ϗ>y�TiK��Jf�2�����
�����9�O\T�o�3�ל���ϕ�'��x�k�.7'��� |���\���<�e���S���R���mZ ��R1�k���m?��ű��B!���$q��@����F�%���:+��<S��H4�T\k�e
=�ȡ}��)gq1���|��Ib��frMp��߾-.���zJ�ʛ�ON��"y]����B��	����'-��l�c�a��8F��������7@k��b߾}8�� G����l�Zk,..���~6.���j5����I:==�w����,i����Z��o~�?������/����X\\��z��%�2,--yd�n��8PTP�'O�G���2/Y���a�Ęh�%X��i,�?�r*C�!MA2zj�sL}At̽�h�ܪx7T򳗦z�kTTǐ&���;�%ק  �4�H#3�P�(�����2���C���i��n��uk��Y"�l;�[0���п�0&�R5-�2�zmχh�ȅ�Ǔ�ܦpF�D,�|G@��#"*���r/��w"9�jԝI�@-����&����uk� 3�m�׫/�̏�׉J�k<�P^����=Y?����=�/_��H	����}:g�L01����O&����i�ih���8���=Z��>Փ̓��ddY���y�|��ظq#|�A��FFF��/B��8#���iq� �}�ѣG155�N�ӏ��k)t;	q��qIDs9>��D�R��|C�C�	�y.� �t��F�y�h?�s��B�T~��{X�����+�"�h����q��|��?��X�|SY�e�崦�|����Y�|D����_�姤Yk+�j<���Q6-�v_٢9�|T�����m\�c�����
Yj�n>���gCs� �u�������n~��P%*�j7g�rR�(��\̑��y�רߥ��4淨Gل*S���"�)�"�	7kB�]�� :���~q���z���Ӱ�4�����a�w���Z��~8Z@]YY �
JZՉ�x: ���E̚�Z��C��D���&���9t�]�7@)�s�u>���J�B�r|�}����Վ�S������~�h[ց�-�q��OR�ڬ,��'�1&s��%���SY��ɽڹ�#��`eQo�P��P����z�����b�i��Mt�������B�UMp��+tS���j���[�2f�SHU�����L�n�/_�%�@��L��B��=L��l��A���|=#��9�*m@&��y�wJd�^ZZ¦M�<�ݶ�g����%tM�#x �T��p��z����}333XXX���fffp��A�z=�رKKKx衇066��l��^Yۏ}��������E��7]i�1>>�n����%/|}�QLOO��h`iiɻ�NNNB)��~�ȕ�8�)K�����0�����IG^Is�n�<����g��-�@xyAJ�>�,���gt� V1"]�[x%�.䇬����Y���L�Z˂��_�/���va�F�I5�w��u�EF�u `��V�H��d�s?�8��4r5c0��A[�jT*�֟�T�ra��A������0�����!&Y���|B�L����چdNJ9���FFF
L��H$tM� F5>>���'����u��n�����Ї>����k_�Z�}����g?�7���8|�0�����=����"n��f��o����=�.�\(����2���q뭷���~7��N���{&DGv�]��_�>���Z�뮻W_}5�������O}�S^ �&-2'q4,MceZd]U�c�x����$��?�ןr�~�z�)�{�Y�e�Y��E�I���l�J��=�fO���K�8ֈkP:V�qnRZ[dY��
��edi�)��N%�, ��
�L��ל :����釈�/Ҏ\��"�WH�@	ZP� ;(u&��TϏ�,�0�YJ!��2B+CU�;d��;��ИT���$ǅ��2AW��S�_�)�gx>t��-4���n�:�l�ܬC�fvvJ)�Z-O#���j��=?�3?�]�v������N:�$�ݻ �n�:�;��M�6��h��)Z�۰a�������;�G��A����i�o��������_�2>������o��y�{���~�םމ��o�IO2��B�[
��}>����a�!n�-i��.%t��	�%��]H�6��O��ƅƄ�C��<Ğ������<IU�#>'��<X�jA�jҚ�w��~;�A��w5�sƯX'���{)h�sD�{�4Ҭ�$s�`ɐt�(˃��X^?b��I�޽S���}{Y������<	��
/9�3|��{2q��~�!�r̲�ׯ�׿�u���o�%�\�׾����o/%�7�L&���w�q^��Wc�ƍ>�rǘ���#�<�?��?þ}����X\\�,//c�֭8�s�1^��!I�����O:���g�Z�o}�[��jذa�_L�����wߍ��;g�uZ�fgg����FFF0>>�K/�sssؽ{7^�W MS���ᢋ.����q�y�y/�f����Xk�l6�7b�a˱�cb|���ZLp:� C�!1u�������Z��υ�T�i )�?p�:?{Zb���M�V��T�s�c�n��Q����)����,�1n� ��S:�6�5C�}�t�9��A�@�>�:Iw�-�n� �w�.����$���=\24��'G�R=�e�L��%����0��D]!����(5��m��'� ggg�}�v<���ŉ'��\'&&�ݛL?�z�VSSS�я~�{� ���k�����[p�]wayy�3}r����sss��btt�v����%�����W\���q���1\}������]<x��z�7Ei�������I�t��W�s��p�9����|&y�������H������ B��7�ߒ6�5���3ܼ"��b�|�	�P;8��|�/��y�u#��G^��)��Gu$3?�3���]��k�2�˴���h�Lf&��t��Fi(5`�n��:��X��Q���"�4͐�
��}�ƩE�t�5�����"�8�ыjP�1�����ɏ��<��8R�Be]�,��\�=�hPr��j��
Z�d�jZ�b��|b�A��k�M(�{J�bb@�'�-)����UO�ӘЛ��"���������S'd��ǕS4�=� �Yi���֭�w�}'�n݊� �������{v�؁��Y��Æp�_��<�9���Ɓ��{�^���<�;�8�����n݊���"�N��Y�aqqѫ닋���jx��8�122R�<��݋f����q�w�}�ǟ6����a||�3qk�_\XX@���w��]dY��=�i�����377�O����SP���p��~�e���Y�\�qp��6^��D{t]��H�+o_��a�yH A�hm���۝�)�&M ۀV5�(�R)D�̎@�q�^���HG�k�� �h�3�n*�Ѭל�y���ư�F�RX� �G0�5!I K��5��Ww4�B=n Q
5?��fL��I��PV�1b�����q�0���x�{I�Λ��"��'�?(��!�7��&��?��x���P���2�&ъ̷�U���B�2��o�ϡ�n�;\:�"|�c��wߍ������7ߌ3�8<� ���099��z�}�k����h6�x�k^��|�#رk'���g���~7�;�<\z�~#����q����SO��_�r�����X(��1�pP:}(v!�(�������͛111���)�z=,--abb��211�$I066��>�����������022�-[���o;Z�j����066�w&���������!Ր	q��1��\*��HXj��ʪ�b9�!g	�B�J�e���B�V�!��.�2�����ހ��>����R����h��W*U4�p��lOZ��ʯ�Z_M��*��`2�J��M��d�p\"T��|e�N��T���Q)��
L�3��	����8ϣ̥����d�e�Yj��ge���$G�!�Y��@���ss-Z>���Yg����,//��N�0��>::�Z����1�?E�$�1��Ů^�{�����(�|�N�e��������;�=�z����������8���p�����|��_ƭ�ފ���}8��q��!��mob"�~��ŧ?�i8p �x�;p��'#MS<��#��������o}+6mڄC��� tp�AJD\�8݄h���2a΅
Ϗ�L�7���*z,{G�k5��$��a�]�
l���i�!�3����b���P�s�1���	ʝ��4����K�P{OZK��o�8��~�� ����@�-��{���C�`S��BHH���)49�JNXn[!��{eB'��%�K!b�z��(")9�B���U�n��vq�E���>���@E��jaÆh4h4x�[ߊ̺�P����!�c=zJ)����|'������Bk���Q:t�ǹ'3�P���B����������׾q���Ƌ.���r�7�_�R}O#Jg�y&�,Æ|	
�655�f�MH|�1�P�UJ�I}�h[>��șL0�,G��l�'�}/\��I���U�� � ���6�2���hc	�h>��)S9T'�z�&�����:ViM�;��P�y�M�hh_%�P��c��Yf�ϡEl���f��,����d.�?D
ƅa��2D<E�!
��2�����cX�U��*=V�)Brһ�(�M�{h���j�:�q�7q����̳���ݻ]���,�'W�q�#sG115�N����y�O�p�Dŏ$���|�#h��8��3q�7�u�{��~�ۿ�~���\s��\v�e��׾�뮻������KKK8p���"j��x���9��a�ı֙ v���e���G������������155�w /,,x���9β?9�����O��2������%q{=7}�=-��! S5d�w߹$_d�#�E��1��V��T���((�!5� �i�����rO�/b�#����'Mk{�/�ت87���=��T( r�(�s'��5Z%/#t��ˈ�"Ɍ���Z*K���H�]�vF�B�����	ג����8
�]H���M�c��/�2.����1ƟzE��q{�y�
�p����t:8餓0;;�ت�\��>B���a<�w*�066�Z���o�?���o�>lٲQayy��[�#Ԟ$	��o�<� .��r�t�Ih�����~����������a�֭XXX�e��]e.��0�"��и�1+�r^T1��V���s���<s�#��M���:�%��3	s�E�\G���z���"q���i��`�ɧ�{����զ5�ӏ�"s��;���s����I�._J�Z(�y��YD��@�7��_��:���b
'i��3c���DX�<ChL�����*��3��$C�k�I�'�2���D.C�!�P�BϴZ-���azz;v���#G<�+� &79
�����ȧ����R>�YE��_� ��2���8�����g>���x��_��=��OŹ��5���1�.����V��W��x�G�m�6<��~,z�&&&����]R_��aii��B�^�җ�3s;��wA��t�z��S
��ҳ˱����җH���w���K5BV�Հ1����ϟ��-?�9�fe�"���Ä��&������Q�6٥��Yk�B��B����L�|��\�|�~�	2=�Al!ԭ�+��3�c$(v8�(�R� J�B9CRh�T!k��<��,��	˼�3�r���U�-T���Fց>�gY_c��EK�x2��*�N1�;����|�b�/�}��#�[b��@��-��׭[������y���jy��()����lق3�8_���}�~��166������_�B������𒗼/~�1;;룀*��U�����' ���'�'�q�X`0�s3j��^-	y��<����,�^��0�ϟ�kRC�4(]�9=�quߩ^am�`���)̸s�u�V;���]"����e�EZ��Y�Z�S�fi���MPk-�� ��9�7p�-��e����� IR���t���Q�꫸
@�5z�.�<)�Q����"C��rRp�%w9^7^'��S��x$��G���c�P��>)l����=$���2{l¼���P�0ɨ�I����n�LB�2�P�d*���\�6��9 �,��F��b���m?Ftl"%)<�(���
����n�q��A,--aaaw�}7���q��!1|j����=�+��W_}���S]h��i\�y���<��^]���$��������@eR?q�#��<�Y>W8q$Nu���t:l7��{�����9(��Xk]TM���$�F�����$��"�4�c��
�r�4Ơ�o��؛�i�����0�S�O)�`��c��Ԧ��}�$�I���]�<#�2X����^��e
�Y/Cz��/�W�-M<e@�Q��d��mYO*��2�H^��zh4�~Oϑ�<1ȱ�1O�n�#}�QC-�,� ��!�M8n���?�Xk�#}��%sﬔ�C=��O?W^y%6l؀4Mq�Wb�֭H�;v��Ν;�H�)lڴ	oy�[�l6�~�zoF�Z�5��[�B��^%M�q���.������$5��l�l#}��s�ߐ�ɵIwUeJZn��	G5&�b(�[�S�t dy����&����c��Ŝ]�0uc��#
���`�P�Hȣ���PQ����5%k�iW
p������!YC�"�f��c��0�j==�kY^��=LV�!�<B������x�5�`֯_�]�3�o�i���-[��t0::�f�	�T!'i���I�.)�=�Pa�p��h4|0�$I�����#�s�N/�N9�#�IOz��XXX�%H8�S��T�ι��P@����@DH��Cv~�\hs��3������*�o�p���T�_�ܫc�OY���B{�B�̟5���,��Q�5E1�<m.�C�J��$2���JkzF������fX;��ƈ�~��@Ff���B����x�9�#8�\�=%}T���Ta�P�D�S񄞗�iX�C���$I!����2�����GA�h6��aNMM!I<��Ø��@��C�����$���`���Z����a$�y��͘���n�����v�������V;v���ؘ?�P>	@6�V�add�F�o#�aÆ�5��7 :��+(�3���y��6����ї���������H�W�����P]ʘ:_j*��J�C�mr>I���4�G`�p�g�7�vKƿ�.���7BX*���_H�}�Ȍ�NQ�>6�5P�~O+�?�����̔B��_�0�>l��E8����!���ԩU���TY�B!�m(3g�֭�馛�;��;��K�7�	G����2ba|��������>����-��������å�^���˿DE����-���(��_}��X^^ƞ={p�-��9�y�����o~/|�q�]w���.^������G?�Q\x��� ��bk-FFFp��!���+�;�8LNN��oƾ}�P���կ~��v~�a���`Ϟ=X^^���ߏ͛7Ck��.P��M�Tqw����u�*j{��ɵ�ؐ��'�1K�+σ�����/{�~�9#�1s�x�LnsU�^�����8��R�)P����u���a>ȵD#�R�t��;�5�Z������cMk���@J�Z���;J����8�����B�\,�y��^]'T�/C�A�tm�&R�F������+�?�����J;({F�i�A��F��h��8��S�+��+سg��%;::�FÝy<==��;��%���̌������'�ƍ1::��}�{���{���v�9�G}_��e��|�_�R
>� ���j���?������`����^���{���?��|�͸��[���w�qn��&��������������H�_���p饗�[n��033�^������B,y��hLңd����2���2�ͯ�F*7gI�Je�(�N7�J����)�	Յח�M�Y���X�}���ǔ��j��X�Z������,�":����,�3�@k(8{=��U�jXC�e mĲ�8�"U6��XU.�C̫E�!��'7$�x>�<3��*M��?\.���[H3�����8r�>����O���F,//{�]�����[�l�E]�={���SOE��7�S��Z���7���h6�����}c������g=�Y~��޽{�m�6���/�S��TLLL��3��UW]�w��Br��C��E�Ղ��N'�p^�W��s�E����_�%�s�9�����8��S���ݵk���}l���Q��e�_��QS�0�_2w��Do�>���$��$H�F�
jv`H��КCHې4I�%ꗌ��~��Y��vgv�y���	���u�ZC[>��LK��ʄ��T��~Ҵ�����T�B�sf�P}��8;�'0�e�*R��9c"���W�'%���a8��P�@�W�GUIN*�B�i�A<�����WY�xߑ���������Ƴ��,�H^86l  |�S��m�݆+��Ozғ����$I�'�'���ǟ��b||q�����_��aǎ��?赉�;wb~~J)�ݻsssظq#�?�x>|J)�w�y�t:��?�Ct�]����̌����?���.���/����68p �Z�~��H���v�:�,�z=�گ� `vv��������cii	�^{-Z������{�v=Ӧg�q�7d��H�� �²�u>�e�BH���5rg���~�F�@��}��\�m˹���yJ�f2�d��5P�$�
Ȟ�%I��8�a�<�9=�h���/����YSW�q6�Z��DP�A=�0q�hd5d�  2)�MPS]��)���1P:C\s�a,�Cf �#�Y�Hi���Uk ��1j��b�.��4���NI��Y���[Z+�t�	�����uN���#=�m�|"�3r;�Д�{ZH����a��1��T�4鷇&�t���`� ���K��\'�r�kz�w��~�︍S�.AT���U�٣G0::���b���lܼ	�:c��g=�Y����GGGq����h��n����e_�G���<�G�sssq=z���[k������Y�a����LEȍuH��ͦ��������
�fW^ye�� ���!S1Q
5A}L�L�(�Q��3D��P"�"�[Ӹ�}��i��)9hܸ���M^�D�7�q����[�����Fi��y��(��#h�'�� cRd����`2Uo!����E4k5�g	�,A1R�B ����8v�)�`�q�aR�D-u�^oq�Is	�h�R�[��$�O��Լ�6pI�o'�.�܀8IE)�|�#6�F��=G�L�Ќrf���$:
��#T�Sz蝐y%D�T/�#��wd�B��d��Żey��A4|-X�PƸȖw�u>�O��/�^�,..6EMMMAk���%"��'I��[��ȑ#�-�V�a~~غu� "�{b*t��1��DSSSx�s��N��C2�����y�~�阙���ڇg�1���v��u����zFk������Q<}b�V+++A�5N+eH_�Z���@�'WW�5M��Kh��I!�b�GH����bi����y?eY��>�~�rJ� ��N�I�;4}��0��#YMn�d6��Ê��OZ��\�u�m]�Pa��Krш�vk
��D�clV$�Т,�o�K'D�J��V;�$��4!U^~B6L��T���*�d\ ��Y����τ�����"-�7�˿������*�F��_�%>��{&��[p��?�s\}�վ����ic�Zgii	 �~�z<���˿�K\~�嘝���FGG�կ~�_~9:��(�����I,//g�4���Y���%B�ܥo��Z�E�>��Չ�'mϼoC��2?�ƇՏ�ع�^5O�ߓ�4Ցǲ���Z�3�-,R(��Y��؞ϫ�C`N�?�AD��9�xӚ���\@�YY2ƸU췁#`�}"y�p�W��w�O�3ON��B6I�Vy_�\��L�L���q��L�v�<�yʼ�s��ʣl2R"������/�ƍ���J��5�W���x�Ӟ�;v�so׭[�������Ғg� 099�7��M �6�MPtn��>��&D�h40==��O>�w�7��m޼'�|2����޹�9�Z-�7::��Q��,�099���%|��ǎ;p��gcÆ�t:~CieQ6鄏�j������ng���� J��Ʌ��a.`�	�*�sNΑ����*��T����)ش��j���ꕦ)b���ְ��l?�JdL�ױ�~�h΃P>ǚ�kp-v�W��}��rN���c0�cqºw�Z����mҎ�24ċ�x@��I!fQ����CV����!� '����Ie� T�C	^'�z��mۆ{�W\qN>�d\v�e�����ﲹ���/~�XYY�\���=z����177��O>�����8���1::��|�3x衇p�g஻��g��(����?��?���{��ӟ�t8p 7�p~�g~�~����p��A��D���S��T<��O�1��z+��ؾ};n��v�ܹZk�}��ؾ};�8�7���޽�����111�Kܸq��]�����?5������kk5�V>_�8����G�C����	�|.2��Y�dN��?�|�"jHp��S�¢�_��P5ı�Tq> P����(�,��8���Jy`<B��X�5ߑkm�h ��*�	oS�a�`�:2�D$��/v��+�����=ɜy]��L����g�БZG���_Hp��e�}�<(����ȑ#~1��x��A3::�wҎ��b���8r���nh��j�|�������׿�]�+Ұ����!����p�w�ꫯ�7��|����W\���;�ć?�a<��C��{������~;�<�C4��	 &&&p����o�6������s���7��k������K/�7܀�|�+x�ހ;����7�������q��㤓N���_�G$��+D|>��+�~hlx��:�n&��r�f\����6���>��k`�s-Z�Gm"t��?����ZȖ��ޣ�
�;y]Qb�
	�as��<9+u��8"���Bf��C��e�<V
�B�c�`��r^?�����ްt���N�̐�Y�AI�m�|��&�d�!ƻ�7(,� ϯ��J�6�4q�u�i6l��O���g?�3�<G����֭[���%l۶��v>��cll��������x����u������a�E���E]�/�[�n�i���`?��`���ذav���w־��ē��d<x��¥��v� >���^�2lٲ�����_�%�y�X�~=����a˖-�����矏�?KKKسg6oތGyI���hx}���ˣ���z6v�hF��H��=��A퀿'=�]#���='�g�\��BE��N��bXZ�5�eB�����H@����Y���*�R��G��}�"�8�y(�����sbp�Ir�PD8�QC�m+��Q�R�1�6�#m�:�"�T�D2A�TU�~�^�;�ߗDH�i2�Õ�Ϩ��ͲL���]�+�Cx���(˗啕����;svrrҟ={�M7�}�{���
�}�ݸ��011�4M=�n4���066�����������{���.�T���9�z��Zcqq۷o���SO= �ݻ����4^�������ή�F��E���z�$��������W�ڻ���-o���" �aKKKx�{ރ�������+��ii?�9��1妕�1u>6ԇ�;��O�	����$ɀk�d�RPH���.<?&��Q�R��Ձ4��mJ!�"(#��|����۔/�4d�b��Z�㠵���P��EZӓ�B.}}a��(޽����gY�8�����8�A/�BC6���8F�5�4E�h`dtI-B/M�*��'n����������Q]�L��Ti���@��h�<O~�/�q�Տ�[N>�����wV�t����3$���Q��}���]�z��݋��qFavv�֭C�������I����~�--�R��seeśhfgg=������{4��Cy���;��.1sii�/��1�ccc��E�5 �5�^��V����"��R�)F�ϸ�d��aR>DT����Z�-�A#�k&�1e�n>�����}��&�uL
�B�C��.��S���q�x.�1�"],�dY�$��|Hg.���*cܹP��4T��DQ�nD��8�]��d6oc�^��f�ܬ����5G�ܼ���\�� ��p-#B����5���-=+��o���o����2/���T��r���o��To��)�$�ݣx���{�n��>2�瞋F��!���C���~�I���s��g�����C����Xk��-BѴ(K§���(�i�V��#G�x7P�P��-..z��C3S� x�I��.��K�I~����l!�<�Z����P6�U�!xH#	�Wv���r�KΗМ�m������,C�[MWY�!�OY_�!���S�T/��:i��Ʌ�1�kҠ$?z�3��6�M �Bi)ԴB=��e�[���WƦCJ�'�n�eDz�l@ey!&�?�&˒��u��c6�Od�!U�,_�OO6x�-{���q��G�v��B--�-//����v�������}��$I�n�:��S����E��@��i�)z���E�NH��566 ^���btt4�^����B>4rl��k��ac��!OH�k�������~`���re�,�,��P���i!��Qh��EPFA�5� �Ⅵp��F�#s��֕������UZ3�/�����U�0x~}q��+�\+(�w��*�d�U�������/{�eHb�ڄ&ߓ�����^�|(Q\{~t_����:�R
KKKޣ����>�JPJ�MN�Z�3w
�f���̌�`�h���1>>�w����bdd�דL
d�'g����4���855�;��A0�֭��t�0�ѩ컜�>��#=]�Id��W&,dݪ�L��V�g�!�\�NH		��᱀xl��`UJy ������z���j��cMk���v�X5������@i �E�Z-B䎲�������F�r���1�2���'�c�!���/�ׁ��R��C�Ieh�wBP��-x{�Z-c�Ʌ�,$�x����O>
SL6�F��(�p����}/�����Ї������wp�e���n�;�����~,//caa�����6l�H���A�$��p�}�ayy_��}ٟ��g��#�`dd���7q�����L����#>�}�c)i��_E�D��=�t� �P]��]��׏��ͼl��� ���+(o��� �8��I�"[� DP*F����E��� �-�B}��"�x,Қ1�*�����X�R'q�Y�G<$��KY�!¡�Uy��<4Cu��ݓ�^N��-KU�jr�՟#�2�Ev����0����/����+��B�BI�(ޞ�n�:������<�������q��<��ø��[�裏zO���������kp��w�^�c۶m~Y)���h`˖-���{�����?��?�;��;��N|�k_��?�������W�������[��|����1.@��oG�Ņ�84�қ-4N!&*���Pe�/��0�/��R Y��P[d�i��'� ��1��.1�Ժ�_��'P�7��Bnk��Z�O':"�l�JVAt�S-`�x8pj��@�T�[h"�I�/.t�	(N8���{�Y^��2�j]+Cs����U0{��D*.�����,��ʊ�M�r�5FFF����O�"�.0�)>~###8z�(���o�SN��^�2t:�Z-�x�8�������۷����͛�{�n�ڵ ��w��w������8EQ����i���Et�]����_�5�r�)زe^�W`�޽h�Zxы^�3�86l��^�'=�I��snn��a��2�nSň�=�n��2PQ9/1�<e9��j���/�˼i\x?��p�*������k]Zǰֹv*�����o

���u�Xŀ� ���JF�3@kd \Ă¼`uȲ���Ik�����
D���BK���pq{�Nc�'�$> !_`�L��a�R�HBD&�1v�L��J�w,V՟������Q^6��4�vx�N~�dV!���:��g���Z��{�����f|�ӟƓ��$w�q����d .��Yg��f����q<��O�&��.�;v���>�)��Mo�#�<���	������o��q��a���ož}�055�K/���v��>|Qazz�]v�������G>�>|����(9��%�ф��\�ʫb�e4[�)˳
��%��S}�[��t��c���K�����DfE�������R��羝ĳx[��.�B;�i͘��o��Z��&�e�u'��4"���zwY�bM#?�V`���XD֩$1 ��	2���.L��2DA#G-n:f�H���=�Cjbd�4TԆ���j��hn�w���^��#d6Ej�����!����iA���(�"'9q夐k$��� �u���RIR]%1J�W�����$�� �'WG��������A!�)r%Š�����{�n��oē��d<����zH�����t:�pn��� �`زe�@T���i�]<x�����,z�y����>�F��#m�u�]���q��!LMM��R�&)��/�т�P�~���yIO���19N�!��\�s��-I��C�����\s �'�K8��9�U
u�i�& RۃRR3�4k �55c��@)k�m �R��,3�Q��������b�&�F�N m`i���#�u@+�6F�-��6"�B� H�e]dɱ3ʬi�Mkma����e~pjJa��'"�2/%qZk�z _��m��?��3NN �h�wEH��e����LY�~(UiE���ǢMIm��\�W�ERS��Bhu�3<��`�����S���&���q���YC1���f�_�'���~��.��ۇ��Q�ر�/$7�ڵSSSعs��<::��g����q�z�X\\�>��{��p�i����Ǐ�c�����h�������HB��e�,9H�R�4<)��x�i�ec˲�9r�e�9XV��^�tt(m�
�����Mn*�~����Mk��ί�4��c�֔�C�ʞ�F���v�) ��YP�X��R�0h�0Ơ�52C��,�q� Vī���\��T�}y�a�&3w5<D ��<^vY���A�E2>[ �>�.�oU����d\$��<�b��g>�Z��7y���4����j5,,,`rri����brrY���l3338묳�����>�{�'�x"v�څ��9_�Z��[n�7�p�oߎ�N;+++����q���O?G��W\��G�╯|%v�܉4M������WVV�bv�OB�[�_<I���8���ɱ+�a�#4oB�H@�AN�P�!���	Q� ӷ�YkarSr=�Q�
�����΃��Z�vf=� k��W_�y���>v�k��	II�қV�F�3rPt�d�
 Hu���9(mz�1��� �bT2I$Ny�ZR���,�/�7H�%i`r��;�I�5(����X6C�1|�5U�3Ճ�;����v111�?��?���$�=�$I033��9q{;-y���v�^|��8묳�m�6(�����z���=�y8p� ���`��G2�Z-t�]�ٳI�`jj
�v�[��ѣx��|����q�	�* �b�ʅ{ޯ�V�L��h'Č%b.c�À�ׅ����� Y'����<�շ_�kg&�uu��"}+�O�/��{"��m>����J�2��V��)\�~��q�8j��xRa=��_s�Ý�e���������������S���~qž-[D���j��c5�n�3��e����NGl��2>�9��B�O�*��2�'��� �8���OMMa׮]PJ��������~����/}�K���1>>�k���zի����k���y�k��»��.<�����|�z=���b~~�O���Y4#?(�"oNNNbݺu���o(���Z�ڵ��v1==���s�:�/��� ~�����c��ѤL��W��WC�ec*�)��a�5L��@�V�Go#_���z�5�a�I�#D�B+$�)(���-Z}|%!H%�;�iM7g�f�������Ui��T�i�/m�R�����J�$�+�wd>U�?,�������V�#���&�
1�P�%�����(b��I���1��^t|b�$>�2i �v��f����`��C�?��w���~���et�]<x�G�=7�|3���/����شi:��$A����͛�կ~W]u��#�����6���p�7�o��o�������5 ����CB3�Bc[�~���$�hE�� }*_z�U��P{yC����	��a����Ԝ�Y�� ��mC�C�˴��XA�12$0i��`�a,��z5�*�`gh #w�R�>���P RXd�ָx���D����j�(%Y�j�jRrN|��D�*��ʲ�Y� T��2���;T7�lB��ub�t��u�1XXX�_�B��%/A����矏��q�q���: �{�n<��OG����M���O|�N����7�,//��j�o}+���155��z��ޓ$����=g�y&N:�$���$�z�3��s�9;v쀵��U��:��']��i����DY�K�#�_�Y��0b��l���1��i�gsA���?��׀C�1�z�"A�v��7}`�u��jQ_��7��~���v�V�j}a�A���UZ�k����w7[�x� �kWHţ�!.�C����J�@^���T�!�	�������.�qDS�;\��e�V�^��������t�C��nOB��nc���ޛg����T���)�z=�i���QLNN�(�+++0�`||�vسg��կ�u�{����btt�_~9��w`ff^x!�(*l����qLMM��?�1��^@:��c�t�e�v��ܓ%4aK�)�y>.��O�5q�`jՋ��1��=�>�\�YCjʄ.��(�T~��yN&Ii���c�֔���H�.�B�ܻ� ��Ъ�����Jd�~�;�A�jw�Af෶��,Ҵ�n7A���Eg㇦�≌oB0!��Qg���P�����'�$Z�`�>'.�,�N��$*����!A>	ɽqP��4��K���@<��d�s�uZ���)���:����@k��5m����z=,,,���)�2�K��4lذ�fӷq||���8|���;�E�>��j��{p�5���D��������rWNZ��'����#B(��O��P��,�'�I�&&��"�>�E9Ǥ��hF�N����dV��Z�s�ʌ���@#K��k�q\�Ȉ�\����wA�ck5g߷Hrg��۵km������(��C ��55���!�
1&�eP��AI� �!
G�@f���M�SX��U*ZkdI�І�v�!e�xCj�T��C����~�U)$
*'{��iI��Bj7��lo��P	&J��)�Ȝ�Z{�m���Ą?4�����F�o#-�B.  F�l6��v��).���{����o�A��X�n���OLL`qqћw�R�����$�d��sd���7�;Nc��C+�'�_h��0����%A�|fؚFH�H�o�a�4ek��=�o�REZ�r�2ШD�B��ϱNk��"�YX���:��!�jPjP���d�i?��ѣ�&}d�A��3e�]N2Q��LH�䌷�B{D���ş	�qI�T6�XTU�$�1�"��D�����MJ�����P@�ec�J!�N�e��\B�4m||�o�j�Z��t:�����;�I-����<&''��-B�I�`yy�fӇ��]��h4�}�v�a��h��D�^�ZȰ�
ix��*.c�|�Bc+�*cR��2aR%�C�m�-%)�`��PJÝuk�ya"X5Lc��4i���1��(@+k�"�*�Kr|���F�r�1g�kj�ᨅ�����'6�C���� ��B�2{�A�H��U�*��P>���G2��~�
�/�B2w9yW�:���e����U�+�����X(�M)���9|���G����#Gp��!�O����$I�����<��}J�P,�f�Y�5c�?��\��[��4J)LLL`ll��B�?�kyy��f��L�~㴵TL���	�i�N�N�廒��(�.�w��%Ϡ��Ԝ9 
	<�i~|��fX�.���z�^U�Ҵ�H�(�dL�3�`2@e1?\�<� G�Z
Yҷ��@�;���?`����2�$�ӌ��2�:d����j�2�:�RNZiK�S^gY����^�!�V?�T�W�?�#�Le��#�^��y����_=���*�{��{�}�v�گ�>��bff��z*>��O��/9�?�||�#A���������v���I�i]�v���'?�I�Z-l߾��z+��g`Ϟ=X\\���~���[n�Yg��]�v����e�<�IOB�Ӂ�֯�	����7�{�qc�e蚏G�qRZ�����դ*���$�;�E���vc���Y�>(Ӆ���fY�4��י����R���JA!
�-��c����b
8VJ�e�F*��om�@f��Cja	����T?%*�B/!��ON���d�����s�/B���a�L>���v�E@Y�2T*��9y~p/���1<�OĶm۰e�l۶��㘜����8���1::
�!l:��Z��F�H�$��F[�n���<���/���.��~����=���`ݺuC����ߎ�����>������/�u�]��Xk}Q��3L�H�Ph��%��5Mk�6�2$]�-VE'!�.�6��P�dY�X��G��|K�	�x��ءv`H��rB��?޴�H�|�]��o��DQJ��N�a��%u�8��F����d
ЮC��A��b�G9�r��q��	-z_�C����O��ʲC�&�@�R���7�lC�ʶ����e����<��n��[��{�ؓ�~nn{�����Dlذ��n��x����}��ߏf����Y�q�غu�_������:99�|�Ɔ𶷽qcrr�_~9��݋x�3�s�=��{�����������W��w�ߌE��rh��s�cΜy�Ps�=l\%��^UUc�S�ƪ��,��F��*�G��$�cG�Ȳ�Zi���	U�7`s^a�4n�������%#��Oӧ˲�I���}"��`mX��[E�ڸm����v�	-�P�D����:@���3:����	�ȹ	��a�:qb		�w�q���~��Y%0B�Ր+C�\�Rhq5�c�lee���<�����GO��E����͛�g�g�ꪫ��׿'�|�g�T&���ď~�#��}��g��rw�؁(���O7�p^��W�iO{N8����!MS��o�&�я~�Z<��Ć�����?? @y�q.K�6e��gC�9ӗ��X�wy
!u^?y����CZ����ס��aQ>iT�s2#G�@+��f��6�Z�cϻt�N+]L��R�%4>�ֵ~���L���fMDY��W9���FS�VSp�E��6��V�5��*t����P� �9[]-#˺���f�2��X��8bc%U���SoL*=�z�"�l!R	�,�!��Sظ�&c�� �_C�k���e�UDG�l�]S�0&�OB�t�bƓ���s��5NLU[kw(]w�~ٞ���d&�փ�˪��O,��R>\��"�K�OZ��I�ѭV��������t����Ą���}�^���|�ALMM!I�v�i��Kp�	'`~~ �I]�-�!�8�S�n�:����j�����w�������%�i���q9r��ߎ�G��.�~�R����$����Z��N��O��~���&@}O�i���~��ӎ�(�P��������*�Tǐ�¯��� �1P�[a/�Ƣg3 _D�հʠެ!��a��*���h���Ŋq��](�C���A�:�ޖ�D��4� ;���r^&���=Q���2�(Cf:�"�:���8�چV� �R��r@�Y�8�K"�$I\h����� �x�r7L����6"I"���#�.v/�p��è�����X��J�_M"�D����p�C��dj<U�[�ǱG� |����Q|�+_�w��\p���~���<��Ŀ�������%��׿�o}�[x�K_�7��MXYYA������7I,mӦM8餓�s�N�Z-��mh���eE8�쳱q�F�ݻ���^t:dY��7╯|�777W(����eA�����#���x��8ݓL�$�Zպ�,�l��įI#�	�T�YQ=>H���!�F&c�100���r�̘�e�7��\��IӚ.��]z>Y�V����?y�u�AC#r������4T�Q��A�:�4B��w��c�8��{���V{S�2���%t�����VŸB�X�-M;�ɿ��y[B�J���CU;�	� 8m��z��̟��ʍ��#�",--ᡇ�M7݄����~;�����⦛n¿�˿ �2�v�m��kp��A��u9rĻ_6�����nc||�Z���H���ԧ������!���q�t�Mx��އ;�������u���W��U�p���������>r'!m�[T�2	�G!���؊C��M�e��T�9!�z��]�e�ܒt��P[�0�{�2S�� � R)��!M;H�`SheP��Zh� XL@J%P*l
 �i�?˴�H���?!��ȓTI��ԐeL�kR�VCG��z�Ӝ�"��9$�`�<���6PƤ$a��}��,��А��5��i��EE�w�VՓ�����J�E�����wm�'��ԧ>�4۳g:�N<�D��u��v���Ÿ���m�6���`ݺu8|�0fff����Z��V����%o0���K.A����� xd���	|�	'�E/z6mڄ��/��L`�$:�z���ߘE1��&0�_�OC}���L��>�i��(5�* �mS�'��_V�)Rk��V�2����h,I���B7{� �&?��58�xdY]�3��֔�s��l�X2K勻.�3# �*��rW��(d��(n *��O��l��\w��Z���w�B); ��U
���T�0\|��D1W��@��«A$�{�Ii�D��-�DUB�l���	1������x��<�X�,Ö-[�l6����;v��{��E�����<6mڄ�{���oė��%<���ǩ��
c�7ǐ�&�e����v����8 ���ؽ{7Z��(��+�p��a����g~�g�o�>�ر��ҥ�@�F���X\\:���VΔ%=�Ʋ�$�q����8VU�� ˔�#������F��"o�B((���L���!C\�H����e�0�E��4 �0fD��z�6Y4��d��;t,Қ�wh�$Y����J�_��Ι�täUw�Z���*���~���x,j�d�:@H���k!b�B=e�����hL�����kY�W˘��4>+++���L������_r&AC1zz���.��.������1sm%I���|��_ŧ>�)$I���i�'�c�����������������f��w
�q��7B)�����ß��������7��q���	h�1???`��ᇐcY?V}� B���X�ܒm��d�C4DB/���;8�z�R���"���R��	͙@ߖ�S5?IZs�%>�B����WE��U&�5��aU��]Y�� ���oj-���Ƞ��٣����Mwݰ$	�����9�z�uͿ*�`��p���������A��u�l���G��U�-[x^ޯb��?��C�r�(Y>�¢'iJi���j��󘙙���}�QLNNbvv���YZZ#Gp�9���(���p��Ao�_^^���ٵZk���*����q�F,,,��[�8���n�:<�	O��ʊ?k~~���X�n��ۇÇczz�{"2'�O�B�^�I�gCt1l����M<����j�l����	N[!A���eD��}>��i��,�E����`�<��E-R�YeS(�@����6s<"0&  ]��{�Ӛo�
�`C%�����@cQAC�����N���|QZ�@�f��1E�}�^2?>al`�K>O��]U��ɉ�7��F�#�~�<q����cٳt�l�A�5�j�T�gdd�W�[n��^z)n��F:toy�[�}�^���O|�s�í�ފ�.�'�t>����mc�E����ؘs�ױ����?###ؿ?���Z4�p�	����?�����p�g������_��_��Oƙg���n�	�ׯ��_�MH���~��1�\# ��YkǄ�;�!.�f"S���3t�#g��E�ǒ$��u�yK�T��<!��P�Da�ud��}��+�
�k-��0���Vʖ�<*�U�[@~j�~�V��Ie�L�A1�5���((�0)m��o�ך�R7��ɠ��b���E�i�,ڽ6T���K�r۠K�6M�?�Q^p���@l�o�0Ɲ�Zu̽D�|rK�h����<\����sXe�41B�i����t�]�'�Q;�In%���C�5�o��<�Ց�'�JcVVVp���c||۷oǖ-[�y�f��ul޼���������1u�\���Z{oҲFFF��t��va��#�<�^��V��;�'�t�1�����?�]wFGGq�g�K_��lق�O>�{�Pb�𭵅�8S1wʋk�r��C�����/��K
ʛo��*��tǯ��C`�v4S]���y��$�U�idp1t�8��j�"�zd��p4a��D�bǈ"@[d@-V0���ع��t�$?4�њ����8ViM�~�^@�����2��WVV�B����|HΎ���c���8xXb����,Tk�̸�Ynڢ2�nG��Dȡ��	�S��뼜2MB^���xVyq��U�@H���%��v��l��EEx�3���ȫ^�*Xk����K/������>_|1��8z���Ff��M������k^�o�?�p�q�ayy�{Q���۷c||/{�˼`���Ɠ��丄��iE�a��+��C�y�����-j����wH0�y��)��q,0C��BTr*�Rs2���6y!b��V���há�;���{�ԠT��"�~�n�7�n��� h��Sl�k������T�,�@��,� ���֚���'�1�bf��z�l^��Ԕ�4^�����P����'��d@����Z�d(<���4E�ZYY��v����Q���m�Z0���Z���L���1�)�Z�����+�d�)-//cÆ ܩW'�p �p�X��`ii	���x���v���燐;13^&�Km���!�����b��]�t��e��gye��Sh��IsŹ���;m��;�R0Y�_q�0��~^/��"�l��h�"jX��@A:�����yy�6?޴��;�+Υ���OJ�j6�^m���~�Zޑe蘗9 �*R��N��D3��Bm�D�=���$�H������vHf.��&�P�UH24�e]龴s�A'c�i���"I���all̟b511c���a�LLL`zzگlܸ+++^�ȺqL�M�����'����I��琠������i���YGjG\��2%M=͝-q�T�c�sB���>e�! $��ǅ��s�<�UVi�y����M2�����q�r�;�L,��A�}'����-'`�v�f]�iP)��PZ#�5(d0F;�O9
�LJg��$�I��L4(!�͉��y�7=O��r���m��@�ΑuY�J���5�i��UU�$r��\ژE'Wi�1::��z_���p��cii	�Z<�O�w��,//���<�M�6aӦM���;155�H�:�	J��kȲ###h����G)�*����z�����^*�:$�!T9�r|��P��������.���
��a ���!�A ��'	�Z�6hR��7��6+K?��}�#�����Z�l�ց<(��2�B��0(�w���ł���'�
��S���X&Tmr�vМ:z���߰gx�x]y�����Hy~U�%d�^-1H�#�)�Gu�W��3�3��B^��C}.�.!l�����|��i�z��z�����������G�O|�PJ᪫���?�q�u�]x��ߍ���8x� �����8fff|����vE����Z#��7�M/���^+ ����I���g��~h\BH��2�eL<��%]�zIz
�U$� 		�Be��7%P��J@���x��
�#���Cs�X�5�,ma � i� k�����ށ�2��Z�,���ʠt�H) S�!WQk�҈�"�$�1@d��0&����q���%B�#�2'���29���6]^?w��Vie�S
+>��B���#�d���ӆPu����g������عs'�?�|oN����M$I�6�~�����F����Z�nB�����y�P|j����χv撀"̈́�@h�ʘ�\'�)��9]��e�\�u���q��B�<�WC+YU�H�q�*���v넬��q�z�-�XOK��� ̀��H�F� :Eͤ 4�,��1, )|D ��65h�*Z~��~�$H�0`�w���u}�]8�fEȌ��S���0�^�����~�}�0�6Յ���݂M��\�^�H(�4fYV�I��H�e�@Y�9�"�������)"q��B��<���x��vCϐi��ʕ�o��E]��ڌ��㮻�wމ={�`���ؽ{�wռ�Kp��a�z�8r�N=�To�/�+����n�c��"��fJ��[&�=�+Z4����*���S��И�gy�^�&��{R@�|$ ���L���|M����i4��3P�����D��/y����CL�X�55�4Gb(�C��`��(�H�A��C�6eX�!�)��c'�me� �a��u�i�^��Y�z������A���`lc#�Z��E�����Ⱥ	Tfaң�e�MDv��D$bu�/>`L�,K@^Fi�+�`!�F�һ��C14,"D
�Y
��аа0i��ׅ����䑥��`�Y���*k�&���_��B�4�����4lf�%)L�!R}Pb�5bA��k��iҤ��NejQ���U�4"��0Y���wl�F���P�4L���|��e�,��&==tW}�J�y����XZ�G{y	��
�A=��o��\���㑇��xc#M?�T�R�n?���ړ�8gB�h�<��y ��Aq����I�dV�d��8s"�G�x@L�3��	���]����(����4��XG�q��:���^1�\�A�4i��c,zP����@�(�M�T��F)�FG�jH��j�%P:�鵑�����z����Ҹ�h��:`���@']�R�$�J�6 ��x���Q	���f�5����DA��I�����8���JA�>��#}�B����1X��'F���i��q�a�J�(���.�G�D��V�� *���B\
,+cX
�I�����eV�A�}~�d�$�6\���t��a�޽���'�)[tȹ�h6���_�e����v���#_f�x�NΤ��'�Q�uކ��C&�X�Y��y�w%ʦ�|3�ji3D���LR�x&�7�O�o!�]�P^�}�D^wq�{��cP�l�;����eT\�b�P���[��"�v=޴�L?M�9��"��i#�L��y�@��m_�6��6�1H�T�qc"��H}R���Ga�����M���Dw�YS�br��s&ƅ��I]��&i��H*SH����Nv�ThHT����oU��,۫�9�ްa����>�s�=��|xc��߸q#6o� ���[q�]w���,lڴ�{�Й�IR���S�Z!d��*�3Đ��'�%/7�7U�H���&$d�	n�' Ӧ��P>���4)�9����^`��㸎(r.�:���{P�ZY!,����.Z Eք�\�i�Jͻ2���Lkjޡ]�@X���H�3����J������Kda�MH�ϙn�����*�ʿ�&�/��&U�<�ah����!c��)�x�w��F�9�e_�Z/���]�I�ԛA|�A<����l���J�0�8ƭ�ފ뮻?�0FFF�h4���|�WۧUcb�\S�&�P߆���A˲x��9>�>���#i�L�V�2pUEce�ED�w�����f�B��}��1�-	�eZS��m��(X��N�����&Y@�Ȝ�%Hm���hu�h�`�J��w�V*�O�7n��-�����B*e�Q��X�<lb��''�<���/'�`ee�&�w�韣�`h��D�1�w����D	d��d���4�Q~}ii	;v����!�"���y�~�E�1�h4���x�3���[�`~~J),..bddd����a�bC�{�#���������#���2��]&�����)�M~�ZY)~�ϕP{=���uun9Ĉ��k�J)�(�S���t���;��ݸ�^��ZkX��Z�������cMk���BQb��@$J��� �s`���|y=�Οy �&T�6�Q����eR���0�G����w9��V�B}υ.ϋ�F�����8}�Q\z��ԧ>�u���<��_w�ux׻ޅ;�7nęg����	,//#���)Y�6W����s!�BƔ$��>��,�j����2ne�.�/e}��2B�x߄�G�Y�����t~�y�8y�<�Cu�ZŷV��%�)�w.g��}cUv����j.���P�0CXkܽ��Y�m(�*���r�P��̸��� ��3Zk��a4;`!r~��VV��Ch=���u��B�Ƒz�>χ3v>qB�zV��ˮ���^��#G�~���� �>p��6]�KN�T��j�	O���i$I���Qo�ٱc�mۆ4M�j�`�E������q��! .�N�݆����_�uZXq��_�oS�� �l\y�!4�Ǆ{�ȱ��d��B48�U�b�,i<�$#俇��e|-ŕ��t���]����`O���2�ª8�"���[�9� 	,bdH�@�+�lp��pk��1Io^�rZƱLk�9�3'�.���G�����9�����DE� �􈑭���I0)�C�3hs��lx+$��}���[վ*�ϑG%�<ܯl��e�*M�P2�2�G�nX!���o|������.��I'��7��M>��=?�1&''�j���~��u�ʯ�
�����h�sr�������t��t011�/�6��5��C�u�}ÿK3O�yR�tB�6$�������)4>$�o��	|A���Y��L˕���\�����5H�Pqa��yVԫ0�R 
!��!7��j�cR��3}�K)K�� ����H�Z2����ː{�� �!� cdiZe�
�Re���Q�s��#�2��d���?k2�|ĭD:���d@��R��2!F,UVb|�V��2(O?���yܛ��ﷁ��9���P�
��M��P�2���K�Z�-ӖB�}U��	�>M�ԟ6533��o������K.�?� �9�?��?�������n�%�\�O�3�袋��<o{�۰w�^���o���둦)������j5���z/� ���]2|�,�|�<$��P��X��;�Q�Ф��Li6��_B�ʲ��?���\
���i���|�y�c���h�����&/����b�Ҿݙ�����:��v㒗W��<O�$I��1t��fm_�,ˀ������	�j �Uh����(o �v�&I�tn>��桕9�J�W�bч�c���M0����1�m����LN�P"�zB�3K�F"0�xx[C�iC}\����ᓡ��P��V��2f]d�Q�:/��.�1�8�����M�6�U�z���'`�q��ȑ#�v�8���166�͛7��3�Ķm�  g�}6�������l6������I߉6\�p�5
���)C̏3��V��]J��$���}��Z�4_Vi�e��Fd�$X��J�H��B��R
�����yp��$	"mЈcĪ�Q-�s�5|��Y���)�+��GY��ڛ�#�򳽏eZ{��kP���*�V�k������se�	Z�����V�r�\ξ�ǨF~�_�jh�P�u�=R�|?�	��BLR����)�j'G��He&p��/G_\��r�$�̢�ᗵ��Od����R�s����͛7�����a%Z��j��G�s�������n���?sss���x�߈��y�H;>>������a��F��u�ԟrU�.RVg^w��%5KɄ�*C��TVg�(�^FSe4���g��H�K��y9��Yp@��X��v�q���/q���2�8^
Q�����H��>�z�k��Y�m����Ak��b�,K�( �.�9ӧ����n[圶h-C��!� `v��=cL���k���$K��v�*F#QZٵ2�B&<ѮJN��V#�e;$����:�Z� ��S��Vfb
����^��`�U�v��q4�k�:�4;���MQ05��엖�<�����������J�!}ٯ�!:�L��g�)	!*�#e��0�"zHؗ�O�<^o���>D+����|R�	���:o;T�	�v��w��f#[+���5�8v&P���$)��}��BB�X�5u�T���r;q=�4
^�_v;�,2(�AY�cm �ǁQN��=t
��D�2DB�;�/]�d>��BB
��z<��QQ9��<�nBEU}Q�ΐ�"�(�9�	�d><r����fff`����֭[�f����I�_��fӟ� ���h�ZPJa�֭���Nccc���@�e�L[�	�2�Zh���k���;Det#�#g����|�׫�C,�2�u�>�����z�0��	ќ4����<�JEH���9}��E��{����QPi�� �ݵ�8���~f@�׵�h�>iͽw � $j�� B�}B#'g�s�9 ��l�%���`����lB�]29 ��Ch����\��P=d��%�C�Q��!�emq{�ĬҔB�T�ǰ�Bl��o�$h6�8t����J�t�I��ƽ�ދ/�w�q<���ٟſ}���駟�/��ظq#6mڄ/}�K8�099��n��린k�.$I�^��m���W��B߫�bDRȕz���B�UE3�����s(T%��?$ e��D\
ͻPx��/>ݓ�Z�h��{:/3MS�j�~���g`p���B:��Lk��e����Gu��|[���ݱ� ����Z���䶳���� !ş�(E�~?�z��1P*CeH)$ddy�l��2f2%�������t����I�)T.�z^2Onk��kp�m�����6>�O�����\w�u���q�UW����#�<�+��_��p�-����=��?�KKK��>���(�9������$�:C�ǪT�_!A ?���¬t^�!5�ZM
�2����#o�!�SU�m�V� ˜"7��{�s�ב�(i@��#0|��q�Q�E��EZ��Y���oEn���Q<�f�dZ�!�� �&;��/���x@����0J� ��/ <���� G�t!f*�]M��5�
�)��L�h]A��+ϟ���:A��h��}/fffk�}����O�K_�R�߿g�}6���7bbb333xի^��;###x�{ߋ;v`������qO��^k��
�sf"�\ �(��C��yɘ)�и����!�zH(��;_<�aI�CY$ç�S� P��5q�m�Z���3�j�u�؉G��ut��������1z?�"�8��lo�_E�@@Ը����~�)�Ȣkڈ:Q��P7- 3�j����T�?޵�ڸM*A\��������q��� �	���(�i�����]e���Ԣ[xAO+hk0�=������۝�6N� m��M�b�@�Dk�#�z= :b ���O��*���¯�)M�Gʓ'�%��
1�'�O6�%����-��'�o[���A�uV�&9ʅ��Z��E�K�i�s���z�񻱰��=O:O����7��M�����N;������_���2��.�<�l���"����_�$Ir{>rW�Zn�q���W^�R���D��2��x�I�DN��x�9�^J�8��L�pp$�Dc-�@���tC�< S�8�h�5��֙B����O���Rʛs�_hd� ���nj�uud0&C7�PZA��X,��ي��6� �3�!0:I�r!�����L3h�N��ZzI:����G��$7aх�5���(����B|�Э���&A�����c�֔�����	����W�����0l�C���)�)x�Z�����<Bxy3���R+���פ�Y���ʥ�}�����y�D֕&\ʫ��.�b�3i�3������|����"N?�t$I�U����V�/�r��r�!�P����iL�������i��T4B���2Z�*[�?l~�y4���`x�ec�4тAhـVB�,�{�dD��\:I�M˴�L`��V}�n�ҽ,Qg�|�(�3�x�3)�j��3eI���1}1�г2���O��ʭʿ������RXT1~�a�x��?Օ	-�(Kʕ��6������;�)�R��u����(���Q���n�}���XYY������0�|���G�E2�2����C�n�ˑ�Q�L9^��!�Q d]��G��p*��*c�R3
�?Tg��� x��:��g�D�� ���SQ5�?���LA�����
����O��)Y����a����$�*�K��9�n�Ǣ��
-8"�V�ʫ�"��򇡨Afb�eτ&5ݗN�U��n�w�Z�r��*��R�Xr���}^ dZ��OM��h��{��_��_a߾}��_�,..�ݹi�˔}JL�3hɀB^Ke̴��|���W���_X�0*{f�(��a��2C��e���n&�1|x�Uپ��{����5.����������vz,Ӛ�l��y�8v�L�U^�<����9C�ʝ��?�v�j��Ys��`��1YfA�t`u謜��.ߑ,�5T	�a�L���ɮf�J�Q�C}(�)���0eu(f�Zy)����z>�QKG)�z=<��ؼy3���δ�m�d#�t���@0���#�N��'����|?�oP��Cu(�]Y^�Y�e}zO>��[/�y�vh��L-���+� s���&�sY�|�GG��y�e��vk-�2�`aimOE�
y��I���C>���6}9�nqCm\�H9fY�6Z� K�S�z��N�I��&���#��:�4���W�WH�����2,h�~����K$%5Yn�6�e��T!e^�<j������ݻ�{��{�~��.�ox���2!>}rd_V.��*A�S��ne�>���ߣy���l��7�<�**Ke�ټM�� ����C�`���"7݄�/[�?Mq̑����;o������yĿ�J�bCI������i�d ,�M�f��Q����"��{I�{T�^�`%��M�цޓ�)4YB��%�&�����'��.sef5}��=����U�w�B֭[������+�č7ވ��Q��Ok D7<?���C2���g��~X{y�K�(g�R�,������_E_��d������v���x�FS�_UP�8pz�u砑;28gǋ�Mπ��[opf�4"k��� �����jҚ2}�D:��¨ &�%���9�֡DB�����D�S� }���%�)+���χF�$��l����{��r�1�2�be�L�R��������&���}��%i�����R�^G��A�����i��BL���3�*�g����[}H�>���0��q6>U�H��qϲ�{Y��U�Ը�+��6�y�9]�|9`�롃��!NJ�y=��c�[=�l�݊���;Z��A�ԵBj2oމ�\��� ��|�z��4W��̣�l~fef�fV��A)�i�������MD,�\�R���(_z�ہy�a5D"z�źP7~ONt���ڔC��Gq��<�9C�G�'y�x��W2 
el�;����[y��V��<n�������o�i���^��|Ozғ0??���Y�t�I8r���?���~:>�`vv��L';>1�4uq���*b�|%�E��;r'(w�u�@�n�J��R�k,7��{!���Yg�ł;b�6 qN6c�t-�_Ys�X�q�=j;?k���o�5t^�4�E� �o�'%�c$����]���
��v���:G�иYdYcj@҅�
ePQ�x^��9��hB��L65�w�����v�Қ"���-ks�� r���\�"��?4Q��y�ΰ��m�{b�I$BH��'�/�I��O��ʐr����F~/T/^F�$!�$Q%�΅Y�	�K�v�j����cFGG��)��ߏ�������q�-���o;~�a�x�x��ކC��s����������>q��n����U�����S��cΡ|�3�q�1���������-���I�K�&/ߕI���{�e^[eu��i+�k����z^�Z-���bcR ��9_�����Q?���Jk���8�m(֎u1�Α�d$���ۦgT&��,�����4��	,j����w�e��fH�q�.�E4B�UF2�C��������3�B6O�/��/�Ư�i�aE�b���s���<��G�6l��^�:�~��>��m�pꩧp��}���Z���	�`�$I�'��5�a� �!�,o7�?��-c�!͇'�`��/���$��T�8}I�tB�)�Tƨ�}>?W�WP��a3#%oΟӪ�∄A�9hL
��q;�x�gsX�A�\K3P�4,"X���tݾ�c�����S�x��@�� ˞��u~�V=3��J�e��!��$=CH��1E�"Ws%�*���UE���Mz^"��@�����aL��~y����*G�C��?ϟ�u�̓3+B]d�XYY���v�܉={��sm_��`aa��v�=�\,--���Ɠ��d,//{dOZX���b�e�Օ�28-H�X���~�Bh�_��r3o[���:t��s. ���V6��責8���q���Ĺ��ϒ��Y?�N�e�l���o�v����3j'�8�ar���3���t:����Zǀ�`"�*�R���|]k�Ydtr�5�~� m3X��C��m�*s�45x�y���LI2LnO��۳9�wi����W��*:�'Le�$)P�U� �(n�"T�T��� p��y������L��nC)�챍��6Z��1h6��@��T%�C���=g���-C��_�$c.�O2l~��["�P>R ��)c�U�L0��P�6������@tk�?.��?�2D���e�?��k���M����6s֍<|��),��u��Rk�.j5[���T���^YZS��t? %�d��1p_�̂&���qoY7���@K�:�f�$��d?�P�@_ޕφ�x���O(�2V&�d*c�ܮZs���t�%��ǵ���x�FJ)t�]_�4�$IP����)M�f�D�����wʐo���;5L������{̈́\G�=��K9.!��Jh�g���M�B��k~��#�%���[I�xA��y���X˾��e����=�~���Ld0�)KA�2��u�x_NB�'-��hJ9;>)U84)C�2��C�
�>aB�PP��L��&@�D�_"=N�Uh�
��R��Bh��	����L�0�g���Ȟ��5R�{��(B�ۅR���{ٿ�Ir�����/���d82?�O���]� �2$�91�2��M6e풦'�~@������oޖЂ6y3��N�!�?�p
�{��;�=�c���z�v;�R�N� K��_S�d���Ȱ|B��ul�Pj6�۠�2�G�l�r�����wᢲʘz�q�{�N�/��`�	��媿�<|!14�o<I����ː�V��XNZ�����T�p�^��F��^��Ol�Z~�6�MD*����ͦ ��r���etM�Bm6Ʋ�BC�1I_U���*˗h�ۮ�;��t_��W-���G�	�6K��u(���۹m�BB���d��c�fH��x�t9J)���U��p��&��@{���Bn}SPY^D/3h4�.�C���6�E�C�&u��[�v�)�.3�$Ebc��Tڦ �)�H��Φ��G��122����F��"��`��~��w��e6,VG�f��u�F���$�P�
� c�uĢt.���iD��4�@w Ȳ�O vЌBm!�#���SX�T�E�?�P���E�	������ȇ�%5^z�7���B���Gc�uw΀��d�u�^/������w/M�E\��=$���rq���W$��0�A���$C��%��̯s��?92�c�+o]�d��ұ!D;��5.�e�8��Xknؒv��T������g��kS#���a��%�+45�̶0�k�k5D&�։\�&kj�:���(F��(��&P��@G0FC�:4di�����fr/�l#u�6�hcy��~Ҵ�L�V��=�s)km�~��	��'N%���o��XB y�q1ϐ�E��\��BQ�}!4*�K�b��~���@�ZԢ���@��89�5��t�
����D��>���u�d_�v�!h�t�3!�(��$T�D� �M��=B�!SH�����%�ʅZ���!:)K��Id^Frn�wCs���'�M�׆Bu(3�zm'G�i�y��s;���G��~ޡ����"ݓ`+�Ǔ�ּ�lz@�(M����_=�U���s�O)D:��
�䮙��|a���ֈT�$5|Ա!�.c~�@C��H��9D�!{�dz��l�e������'z(#�P���B�@?ҧ��!ab>����#��CcjS��a�?$��ˤI�B��<C�ec�Wh�d�<���Q�@�3�P�qZ��F���B�����x��1��֏�,�`�qA�tq�3뀜��>!b���4�IR(c�-�-�̱����g�Jf��EL�Z�B0tla�����PZ0q'� j-Q�9�>�B̟�v�ȫ&[�hmQ(�����MM��x]��xH����:�6V%��*�Q��Cm���		P�Q �ȮLh���)����W��6�w�	7n�!&���I&)��0!��e�4t�R�	�� ���� �s��2�4�c�:��?����)/<�?�T.�z�0p�X�oΊ�нE�\<}�OEm�2�CR������5�~"�5�զ��[�sbP��Jrb� ���/K|�Bv���C��q�C�!�
1��Ph�J(��Bв�e����.�p$�哋/�1�*A*�>�r�{Dk�߈醄�*�@��a�/�Aٶ2:
��|V�c�����Q& �^��+������(Xeݺ�.��&��3ա�(r���$A5�^��\�yK03)��~$��/���5e��F�!sw��`�)M����in��]/1ŝj�Qd��I�	�lb���T�[��(#N~���P�Ԣ���=�i�G��&T���Bm��ч��j�VC�͟	����|�v�ߓ�������x�YVY�b��.d^�4E��7��B}�	>~�_�u����KH��C4Q���Y��i!�V���6�)�{�6p�%���Ǔ�<C���He]<}(:I�HTJ���G��h���0��M�����u�`�ǳVa�����U�B"O~�ɼ���9�����D{e�CnÈ�R��!�*��R}�Hٗ!�!��cD��tM�4-C��r��bƜ��{4�C�G��Cڹ����u��i�^������ai�!b8�S�I�X&���e�B�c���Z�N��u��u]|�y�9�����A-��ę4�]��`�^�s4lfa)^�r�f��]�u�J�B\+�x�iM�>IW�� 	�E�|5۹���VRGS*�1�L���{��2OOR���=���'n�$U��b�!�%�Yۏ�M�3~��+�!�/T���0fW&89ӕ���
���"�MY"����3�����e���7�b�!�(�0o7�O� KfY~������R*�TB�Ke���K/Q.0�A��CW���%�5�b�r��V.d;�廾�F�F��z��?��^(������/S_��@oZ�x� ����R@G�����A�Q�)�$u��-5�4�ln�I�招�3��$�1���Y.�#�a��Z���JZ�w��:�#��拧�Q��i�;�c�7C���EH�33���qN�J�M`<�|H��a�=+m�?�%��d�%#0@L�6� �p�<� ]����%�E���B�݉�����<� x"���Iʃdq�G��>�چ4��߼�!����
�7
?!i]�5^x
9<�J!.�/W�_h��?n��2�(�������t�燂���X��T�4�@��u��0�Y c2��s��h@�2W9X�AY�ָ͂Zk�� KRhX(k��Rh(�h��y�i͙~���yp�K��E������WJ��H|��!�Xy�b	Q|A����aȈ?�30yC�j��+IA�F��VnU{����BY�P�ƃ�Q{�!}i���P>F\���#]��S��I�7�Gb�$�Bk.��dh,�P��������F�ɀ?���:��5��e�$���U�Iփ�_͚Oek/�9���vx�3�%�:�h�Kh킮Y��������A��Ǔ��e���0B��A��H�sY��i��")�OJk�����E>L����D�Kh(�!59� �G��?�Hd!�^�'�dl�{�I1�!P�I�r�kF���c!��2�Q�{���y�P?�ߨ�ϲ��h?%?���.�,�����Ɨם�+ߧ1!��`����� E�K�\�)�l΄0��_F�!p&��Lg��e�e`e�oه��}r��j�:�`F)k���UP*��	�j5礒�
Q����FŠ��|Eye3t��R�}Z�7���i�C+ї�(r-��+&AY�<���pX��Q��P�5D:�-a�<~-d���c:.�$�|W��BFe�J2���8�	�ći��d��~)sw��rX{��Rʫ愨x06^fc��/��ꃲ6�����xs��m0Y��e�BB����լ���Ucʟ�m��s�|��B�O�b��>P�m
��5�6ƅAQ;��,zT���X��������@f����Q�D�|g�N�����&��Uk�ǈc��\=G���ȡ|f�(nq.C��h��C��U�>��g!�^;�G��|�j�@�L���e�7�4���l!��yP��@C�P��Ʋ��1���2Bm1?ʇ�+�~��D.�̒�I�,�6$PH��~��*���B����#�'��*���c(U��%Ɔ�{P�>!X ����Y�]Xk��<%C�k}��wf!�0ơ{�A���i���qgG���Đ3��Ike3�^�F��K����ɾ���C�<�*tk�b�>��^�I�:��441�o=8aBȊ#�[&^7>)d�Uϣ��gy�ʘ�|^^�Q�Cɔ� ������zq�>|qV���Zf���烬�����P�0��ߓep7W�,_')����Z���m2�����O�N�'�;/����A�4`���8+̝��e&<ǉn��X�����laJi=�Ł��ȏ!h�9� #&��!�7I��ym`Uqr���Pm��y���=��c�u�v�1^�� ���K!1X�`��9s�����P�����0�.�G������M��2�&�Ƶ4k�?��/��ze���`�h}��Ia.=sBBZ
�2z�b�e)D��neu�$=�B����;R�P~^�1��L~Ʒ�5h���E����X[�v��*�G
ڟ�{lҚ�";�@<���w?��z}�#%.�hq�ޓ�<�
?�ʓ���˺�I��hsȾbB2�2o�:��j�M����sÄg�����P�M��y�~��zZ�vkYN+�L�v���Eΐ`�k��;.�x��8F�V+h��I��v�1ei������+Bf�*:��Bh|�Ƨ*�ƅ�cY�H�Q?�4��\՟<�.�_�^w���@�߸�uy=$�����5E�Y���TTG\� 5z�:F�id�%D�:l���X ��#�]05k�Z�T��2he k��d�uX��E� dl����P�灊t�QPz(S����_��Q�)RS�\�B׸}�>\���2fv�9�b��I)���k=$��}��:�>I��r�!�B#܄AI��Q��5�Y_�\��G�^R�S$�,���с8yԢ&�o.�T1�<���E�	��/+��3oI��k���~�v�u[.nJ�|9�y�ttcE���N�306��Z~�*���PF`���4��6d"��! �~�IS�=d�/��������].(�_
?z��7����4�8z�����X@+��0vs0?rs�� F\w�w�u��Hk5d*Cͨ�֡l[WH���A �A�)G��,t0��:+G�]i#V�$���0=��q��_��4�"�-l�����U�B8pB6���L����B�q�o(,��Ќ �ְ"n�d�2���j�/S[B��&G����̻*I����τ��)\�oqRzw��e����YG2By�5^�g�1.�9��em��"�	ч�лU�T~�c�-YO��0Mo��S
�=$ly��ɾ��e;���O >`aU�ZCy�>دQ�"|Fv1�bl�AY瀡��i�/�)x\�E\`�����b5�6��q�"���7(�k'�8i�L]�'�h��l�d�!��!B�eBBj!f[%4By�ޫzF�W�����)T��_�B�LXITI�̎/ߕ�^?$`	�s�o5I�� I$�6�.o��^E;!�1L��U�챤��T=���2R�>�@���e���췵.|�����:r��r �h��,�[ˌrh�,���(�J���iڃ�Տ(��O�y�o����!�� �] @���Ţ���F�^G�1V�X�}�� �`��A�$�D&Ɉ�=zg��,�+�)�[M]V�7}�?،��m�����_N�P$j/�O��!x
���Dsd^�&@�'i^�h��-�(S��=G�a'����ߥ�����V�=e�X6_�X����2�݆�|���Z��4��>A_˭�4"��i3��*����A4<������_�V�����۰��DB�ӡ�A���&I����M�q�6P'�����6g�\���b�;�M�Ҕ�Ӡ��^����u~<i��Pk�d�f,UB�M��=����>�̏׃�P��� ��4�I�q1�a�.��|O�`����{��j����j��	��	E�7�@�?���!uf�49��[��&���R�ݮy��;�R��4(��RQ�`��Y��,�6���"�3�'M�%6��"B,y⎔�n"��H�>�Cy{,V�e^B[kő���|�!wP�$Q���[�lK���eU����rN��י��x�36��X�`l!Y�,!a[���3 �X$�Ń-!��26�@�YHH� �۴m<�==���ݧO�۾�U��2���X+VT�����C����W�ʕy��222R�nm�I^/��"KP\����ք��]�5�Q�`?w��9ެt/#p���+��,�9(�v���������h��,c��gz����R����2_�6�D�[y��]��_����Fe^���rX6�ϧ�>x|�xAJ)�[A-.+W95�uY;��v�OD�&����z�dYt��2��6�I��q�2RΈ��!�����j#s���X�T\�9Ax�����qV\O�����U�5��<,Aޚ��K��i�]>�����@��R\L�K�.�@Z�����A+��g=o��|��z��4���|V�}��X�M�����P�i�YϬ�s9�_nsX�Y;��Ap�M6}���9#r��	L���eQJ(��r�#��J�;�h@�Χr��V�WAoT�U�rG�,I�_���.m�c�߬����E�֥t()%$_B�^BkʡUo����,W5~�;���5ZCu�z�)�5.� �Ƨ�^O�o�ɖ@[S����ݝ���O�_�!0��D�-;}Kȶ��l_�([&>����I-���:KAj��(͗^�H�-�U��h��y�JX{ɱ��;�����5�6�q�^x����I�x��rq�F�ODŻ�A�d��>wB�=jhr��5ܘ�j�r�obԓl��_���x�K5���,}���*B���__��lp{w��G�ô' `�q��I��%�x";��55��28�o	|�+Ѩe�`��u��i$m���ly�A����fo�w�=,�''�|��3h#__j#}ۥ��JX�ʮ������ː!�a~�e�28�m���M�uQ�T6�O9�lm��w����o̙Ӎb�ȶ�B[���E�?�������<�q%��q��!Hc�S@=9��*N˼�8u�R�Ki
�HDp�s�oj���q��}���%�4  #v ��Iٗ��c\� bٛ�{#^�1��'4P���T �����u2��C�?MJ�<��'c��7/.� O�R8I�!]9��`�����<�t����f񤑝F�9iS���Zd!Q�R�I[�f��!h!�5>���E��5���P���^򳖏���݊=%ߑ���������U����ej$�O���o�����[y��#��go�k��r���6�V9r�(��P��(�T7rK{r.W$�k;�濛l�܏Zu�~Vz�BߡĻ�B;; 5�Ir'���F��#(R9�X':��'J�Ƀ��C9,�RF����@ �z伫��RhAcMF�*���X��<��ҿ�2��r�*Q�5$���n8U �o�@$ʵ���OV���%�[�W
R]��%z���O��v�n��?]��J�}%�O�����d�uZMk���ZP�H�+�kޜS3p;5?�����c�9P{~�YE����|S�1xTA.ӹ�\�U0�Q \���	�Ů?"�X�����st]�&�yg�������@d����$�i��|*�+��c>N��@���%r�Z��4Zj����Ia�BeS�a}bI�[���-��D��-��ٚ�-�"?[
f�9��#W�f�.˷L���2�I���v�
�%�ׄ��\.{JY�\���h�$�^2�-SY�,�k����D̍6֦'�/�������?�|:�����S��?Pn�r��?�e6�^�})�րk��6{��9�E ˃;��s@�hӷ)鎲������R����Vɍ4����z�Ic!`kжx�F���J#�b+���2�}X��u�����/��yl]�n�w�m����k�A*�]=&�s	�sZ�WJ��-�k�A�o��'?�������Si��5&Z�  ��%�}"�r�� 9�\���(��A%����i,���=B�����e�#���[Ɣ�DT����,��'mD9O�1r�H�4 w�Ь;���'&c��\	k��4������2?�W"�K��Fg2?�{��<-�z�b�&�����5a4:�N��9����s���s���ƺΒɃe�רQ�d�Y�����D��-�;�����u>�Pd�H>u豸Zʄ�[��5/ZuӼ��F'c�-���y�[��0��&�rdT`~%/+��#�������f�v,�'�� �Ҿ�S`�.'���.�Q��<�`#{o����xN�^"�-D���S�у�T�� ^�M]�WK`�i	~K�Y<J�<�ZHL#�K:g�k�V"d�"�#��_-!���K�%<���Щ�^�<JС=`d=���Ɔ�&-E�}a�n���֘�f9��l�	9��}���}�����G@FB�<�������&0��?y�zs׫�7㧯o��s>10���Yx��J��Fˠ�!���2�3�b��9g����a�ɖ���.�pbg��JC��Y^ �}zV����9� ��Y H�$���xX<��{��΅�<�)ZI��D�����$Os�=>-�ۆI����s��v������T�%���/g�?��Z{ZJ[��$]-hur�A��7���+�@˚��x��Lﮘ�Y�O�9��:�da:K����_q�ʦ��6�{��{sV,��\��!t#��ؕ�=m�; .���:$J�-  �y n���GB�{����8P��1�2��iD�M���RNp�������k� �.�X��'��'/'�\BsY\/��RB�X$��N
�j�)�����Ex�1�_�ATVv�y�x/�� ԓ�5�'���rncR��m}�x�S�B������D��sd۳��f�Y��3�����D`��s���>2vOZ}#"���}w�'�RI8��7W
Ix�e�q`�|oC%n�q'>-4/��x�������y���z��V
��M#@��|i��J������rgv��Z��{i[�)������v�Ҙp���x�p|��� J	!ށ�C#��C?й>?@Į���m�>�wC�r��H�����!g�p��bXB/K�U�k{ݤ�A�Δ4���'�V�-��ZSk��%i!��e��,D!��9�P���\����Zh���S*6.G����Z��Bƺ��v��|����m���n5_���
��{�u���Ku�i����\�EV6/��ϕ��S��vy��[
|ݮ���cc)I���<V�ŌXM�b���N�dr=��\�+P9J ����,�9�����	e9'*x�������s?�4��+��TD��������3���ܺ��s�����Z(���k	[�.C#-��o�/���S��5��-�D�#��)�5�`���\֘�u��|.WW:�,C��j-@YHɶ���JI�pn˱n�rN [�,��(�Q��ʪR�cDpK��R1��ˇeK-	p���W��DF �y�k|~��������M���jN<;C���9�9�l��˦����x�����Mky�ʇ�I;mK���yn��qٖ�Z"#Y�O!I8�PZ.���YJ�j;��d	*�Y
o˥�,��?���V*]͇,K��������ּh)�KI�סd�js[�����M����?�U��+�l�c~=�i��#�He� ʳ�cf�S��e�
}6��A�ir�<�nZ�(�t�B���#U���� ��nTk��J�C�[�˚��[
�R��B��bkRZ�^nlZBcM�97�T�R��%��VN��ōl?�J�x������BCE��%i�`���)i�yhd-˵�~�gk,I~�<Y���Ĺ1#�Ҵz4�Z�K�[y� �<�rt��x�H�q1V�2�:�P�אַ  � O@Nc�_������A�U�r�^
�^�^��! ;7	��y!�)S	3
T���D ��R��w�l�ĒZ�;$醽d9uN0�3��_�ZHV�'7�,�V꜏��Z
c�a�K�v�nk|�޷xZC���_V�5�$�Z
B�@K�/�G��P�uj�ުcK�X}���t��=���������R�\��%�l]?y8K��;lM���\��M	���ཇS+��\�j鵛w���;Uӎ/q�����ӕ���F5J5r�R�D���\�4���N��d��\�R��;��KӋ�׃C/E9+��$=�4��]��=��+��ʱ��e���;:_��/�tJ	>�]�Z���yYJ�B��/���y�嶔�/��|Ƥ�{-�l�彯7�A���H�wd��͏�@��ܖڛ�9�@���Q�-H6�M��"�#%�6t�+OQ?��R�B��M[y	}z#~�Rs���K��ݿ��:P�H����ܜ~M�/�����w�^?����,�"��tK<��-Ac!]�,y(e��C�/]PY�s(�54g����,���}\*3]��ޙ��ǜ���%�t:����4���,h��eV�K�`����( �����a[|Xe\"CZJk�:_w:ep=��w]WCo�q���#|���l"�lw亜Q�,L��}n�>O���v�#�)1�O|_ms)���nH ��y�u��-���؏Hi�]PR��v. ��q��l"(s���0�=����ȹ(z�k�����u���].�@ba�.m�\ɗ��>�dMkp�I��0����Debӆ����L����4��8�ڤwI�[ʸ�
�d/F��~gBѵ^�s�>����??�}��I�>]�y^�� �J� �R�̀2���R`�g;xl{�1�tB�٦2�0��������s�<y�*��l#6�����(�;
B�Ĳ^�)�D��ˤԼ��#�K������r.��A������ΑHR�� �XC*����q�{и�Ay��Ic��\#h+�ز�4r�d��B4�.�Z:�-��n{�
�eɺ�x�����e����~k�^�����n)=��=y��Bu)��m �VƒO;�S`��	��5H���?�����H��F�2�>ȥ��qǭ��g����X�q����OBX��ۧK{�O+�b
�����fK>9/���=��WI��{�%� �!S��g�_{� �i)�T�=@�#��3~�
ɉ�	�ө�!���Y��ֈ�IHFL�4���$��m�%�Z��v�_��HR�(�q`�R|���J�����bhO�ӍN�<uR�9wYh�E��g��e����=��$�׊���K�$�>�M�K乶�x?<�|�nZ�j�sL����#�b�/��c��t罟OUك,�����*�l�����BV��$�:x�ŠL�_U~�
���@����-��i��-�6!e���.�U�D^Fi�H�����^�ٚ��5�,����/CV=$i$����|-!�7��l�����п��%du�ڴ�y��W��v����g�2�<J^'>��\����̅	��L �D�|5���"��E:'b�aE�|�q*�#}`n��*�G��q�]��lئQ��
��n*'x��?u_���"a@��a2,�!�ք���zWO>k���?G�ׂ�\~�ri!�-��:����XC�-�9�K�rM��|ZB��j	)���B�5��6_�kJs��ض�����f�t���m�6��X�iel)N#W/��C��7/�xu%�o��1�P��}DJ���v�Q��,�).x�B_�ύ�_p':�V0��z��U�!���% �l6e�Ѽ��f�a���Į���P�i4�\C�Қ�>�D-�������.K��Ky�Э.�B�-�i�KKH�[EX:g{\qz�DO�)
�i�f��~�2���[��2��a$�֟z����3��U��S����?.��X����I�Tq?�I��r�k.ᯓ^��Yo����[� ��m��������r	R�^}��s])B���ը�I\BJ�;��l	�5��Nv��h�#-�=��d:-X���h�:Y���->[i$i�qn�[��a�<���1�T+�^F	�6����|��ŏ?��=c4z���&�n3����Lk���V]���n+���T��Q�Yk���6Wɼ,@�7�[e�vq(w�G�Y�x��K�����Vk��R��2�ڽw,��i)s�:�9 Α��V;G�L}�)�P���� �!:�t���-�*�뉹61�3n��l�V�`���j!��-� �yZӵx��Y�w��L�_�qI�kMZ0iZ�'�@�Y~�x��.��˴��Y���e�i��kktne ��y�q$W�VZKXJ��Yͪ��-���i�R�wU���ß���m��K�5?��^��Y1���\��H{P�Ub��y 0.Á�||FNG�@��R��v�c,��o�w�=R��#���k ����=��A�E�m��[16���җZ�veD }�٣AOP�t�w9�� e�������S~�M��G�K�2�+6���\NIk0��,!���n�<�*�粟�Y 釮�nJ	�);|]z��R�N^K��:rfaP�_΀s1�/n�wj�ў2DT��F�t�3$�%�=�rӀ�i�zq���q�\9�����6�� �ț�׾��m�#�0߻�4��|���MsQ���B@������ �s(�]����4�@H��p��'��P��сRB�>�t(�-\���-��@���k�ȡG��-�z��
>��R��� w zs5�p�q Bܜ�駥7������O�Z��Ϊ�ܩ9g�X:��:�\cF�p��
��k����@פ��z0Z�]�#��������B�S۝��'�u��ߵ�|ů�=)5ŏ�&kh���,�P�����g��x,��(^
�KP��2���Z�/�@t�F���G�O=~�q'��5^t>k��{�`y0���˹�_c�S��zo����ri��xb��Ӌx܉�:�߹�ק�7 �'�U��ߢ�)�rPn�GFi�P�n�/7�;��!��ExGH�8O>Wl�ι�m�&���_�$\	!:Poo$��%��t��A�?[i,a����?[e���ZIX�G�v�B�H_�&/����[�[�\~��ZJ�RnVk�h�_����T ���e�ւ���|=6-�� +��9�ǡ�{N�[�I�JT���wI�_�˙|��@i֬�s��"�N�SJ	>̠v��̂Q�yF5Jd�W)�_���Z߳���h Wla�v��oز �G�ID�x"p��S�{��J���%�Z��B�km�y�b�y�r�l�~Isz��}�����ZK��Z���e�d���6n�MkL���"����%���^q��[<J�� ���%�]��k�����7ֵ���v2y�C%p}�ˠ<�� w�S��.���rFJ#6qi�X�C�u�U�'�n)��J���T"f�v��
|��\�z�b=��|���\ 2y�D rp�	�;��G���P/���y`��.�A�P�J3��P�ʹInLID�=���Fx����<'���[�k�jev�Q�s��:���-e�B�k�[nkH�'��fE�nzk�k}�~��A�{�\]�jo��ZHY��H���V�5@�d���^�r{���?O����E=2�1��,�D�sh���JO ���k��e9-�楡.^�^�ЗQ��x�pX�!F�����a�e*��JP"GW:+���1-P¥��J��`Ԩ�����5���]2��wl$va��,�Z+	��_��߉hq�_-T-��!%�3B�P����������W�ǜ�U��Ν�д���7�����ޥ�&�-p�z�?���8�%�:���qDXU�q�u�R�;�ꢡ�؅lP�\��b�'7�z���.����w�.'�)����Kp���@T���5�C(�����ȍp�Qq�ʳ�ǣ(��"B�Hc��.����/Oд��֨���-e�'���Qڹ�d��gY��c�Ё��N2�|=x'���su?���D�J`�����|[�;7�D��m!ܵtVh�V������'�����%��%�-�t�=��6��	�UHpK��b�ճ�]Z�M�8��O]V�$�K�e�x7{τ�itY��5��y.sG	a/���@!��L[���H<}�T�Շ3�W�������&o���@ʈ1"�!�G�H�)�a��������%t^��Z�]2�%?Zi�!�s�[�T����������Z�[[\��Q�U�r���rX��h���J�P���)]ys����R���$���&�t3��V8Vޖ2� �ڻ�okʗI�5���z�7֪��W�kE�\q{�9��ѣ�o��;d�(��OH�a���6T��b������'*
��������.��~�Cؠ�޼�� s�$*����b3��0f?�=� "l�;o���1�?��p�tb	777؏�At�]�a��C�(����J;�*�c����Y^��$�h�ޚlrP��[��%x���I!,W����,P�]�-N�jĮە�Jtz0H։m����̛#KZ(�%t�s�����e��J��`%/2���%�%�k����"��޸�1N�����N"��Z�8��U����l7�w%��K�ȶL|z<�v֊�,�.`�D	��(c{t��c�ǻ1"�M[<��@�MG8O���tf#��H%tD.Q��].6F����=���C�yL=^�Q��F|Lι	�/&+�},��5l�$�P�l6��]��C���["�V��L�a���BO�5d��-���C�(�YK�Z$�����K��Pj�}k��oIY����$��O��o�)�Z��k�s�z�������%��.���Q�����N�ǭ1MTLz.r=ε�ڪ��ߢ���4#n�-�uR�f�� B�|�8�9Q۠2a����Y���w��r!0h�l �����A ��ڪ�~���ƈ�Nzш���wHc��w��T�Q��)�n�5aku@Kh�/WZ�hT'�����½%�K3ۉX��ˬt1�7cq~V�ɉ���+�ۦE���лt��Hk� .���n)�yWƸ��^��5�d��K�J�ZB_���.����Vr-�֚#�k�����!�z�����-�d�c�{�\c�O�W�O�>2�,2䰼8%�NȀ�����Y�,�v���K�X�<�1��`�п::B�s�4kЈ9���x,1I���hX��P�V�{�v�k pk��g���ʰxZC���|� ��V,�������<-����N�\�qN�S�kB�����ZhVn��Ƨ�vZ�a,d_�%=��V�Y�Xc_�#���Z��5[|:W+J����6�� ,�w�:L�N8�sQ�B)��,T�+�sJ\�T ���n����WA����ʼ�H�-�f�X�a
����i�3#�a��H��qJ	c.wnn\����r��*��d&�B�-T/���5�����	9�X��m]��
A��R��܅P{Z��	�5e-'M��)-�>{Ej	9,��R$���x�y{N�s9_N�ɹ����-����V�Cx�Ϣt4�t��}n�Ί[������r�/����e ��U	��#�@�^��\�P��s�p�N�����l�:r;�//Co��܅�+˧UML4����$"��ݔ��(!�b���=(�i�|�;K�T=)$�rY�Ū�%��P����&,e`��F����,����=��f���J���D �W:�U�V;,x8wG�"��s��R�7�ܪ;p0Nz��O���Vi��1�R4R�ZudA%�4��.U��E;4H�9��핪s�Bc��R�z���(�yOs���t�� ���)���P�B�:z�B?8_|qy�-6 ���\��g�s�T\��g		ٕ�	�U��qFZ4M����\R�kD�i�=���MI�ɯ=A�������,�4�b-)Z�R>_S 9��Yk��~K����xߪ��vK�a�0��<��0��J�R�V\��f�Tڥ��X���&�u�,~t���ksM��D�k�@�}:Nئ^ۆA&�ˁ���]�y�&d�K�j����ؕ�f�v�8�9����Jo,���,��Q�{1冭�W�%T,�����9�=�P�ʺ������K�H�0��К�	�,�x��Y�k>v��B%�h��5>d�^��s�+�hKX����[�[����Yk���i]����6���.�(���v���]kE֫ՆZ�O��7�-�5�!ؗ�r-x�ج���S���\qI�)�|�/|^�wo�arcs����=M�+�,���N	�;�������.��.���G
��w � wW6k��@	�� 8`�����mN����-���:�L@ppc��2��Jæ�w��mF80z��E�r��}�C��rG����X��/w��ԖH_//����-�`�AY/^rr�(o}�N���\��l0�̿�z']?3����/
�>�wyɫQ�#�ĭ���k�yՎ�?�m�Ֆ;�T��6��dk�F��^�= �_���b�����b���i����-��x�V"�y��/��*�S
z)�=�rk�rZNC3��=:� dpF9J��
_�X��Xi�B	�t����8r�Ā@L���ץ=3!SB�t�� �#R�i�+zP�������c@�ẏ��3t> �F�ܣ�!wxU�F���?x2#�c��Zē�{�<��~/'��˓�ӠJ�~��S毑�$��ɯ��Z��B�:�h�Z�g�u~*�@��V�uy���
 &�C��,Ī�g���]�Y�5=W�hem�!ӥ3^��X}���ƞ._��9��[���r����]�;?=�O��xߚo�nU��O���z�6g���j}w�z��rק�%��!�/3o)%l�F�,��I�/A�u����?����1�K�qDF �n�'W���$�	��U�Ý�vq�@DT�-��@ 0���mL�g� "Ń���]ݡJ����v���ޟ*��4�:Xu}Y�yh������y���w��s�\
�`X�z\]"�o��s�V��������&Z�q	���i��Χu���M�_������\Dq	(�>�˚\�@_ˍ5�q�7F�8)MDs`?G�P�tV����*r����<!;Bv��8>-�v���l�MW��D�L>����g��b�cyB4��l+[^g� ��A	�5j!-�\",�F�&�ѓ���J�Fx���CNXk�Y�ת�&Y�KN4[vZ�>RIIt'۶%�Z�F�p	i����<�Chk���D!YyX���Q�����KQr�X���r^�k�-�Y�ʹw��Gk|\R��.Y���Փ��rK0!yX�[Q�K�-@J)�բ|���lz�8��^��v�d2�~� P/4��2<r�����3�Hl�v���pu��n�a��#8��Z`F'.������Z������o�vsk	|�]SkR�����Γ�tu��$���H����Z�/ӆn>q�󐫯V;X��Z�j���&�Zk�KS����jg�?Z��V�-����{�}���%ح�����V�h�d9z�i�5o|�d)KM9I�O�z��:�E8t�H ����>�^ B	�� �9�6% �"�\.�5�*�4�+s"� � �?g�n�#�|B�;�B�F f���-(<�^�N�2K.��&�&�XZ��ǥ��R>ZI��XIz�U#����.������zsO�Y����b�P�nc�2��Z.���(�V�O��NWRk����xk�[e��#��ɼZ�eZk�ho��2�w�0�x��ɠ`����.���������r>�+.��H�����\�"̡���\�6�;�\����y���7Z�t�z�E�bW�a���LS��A>���.�i@Ln��c���᪞ƅC�4�U�.%�֐��UL<H�qI{��.�8�@������*1k�"�A���a�$���7?�vZ��5�[&&�LX
k�w�o��%d�4�Ч�������JAo��gLZ�[cEzk���4�i�
O��4-e�ǣ��E�`�Qyv]�ח���r��}�>8Dko'���I޹\ 8dG ����%�&/.��*�x�H�]���y��e@�=��=<���6�%��a>A�@v��p<Aյ�{_�:��ڏ5ε�%ۂ��Z�[�,����.� %�$~Y�?7�,@���_�ҵ�p4b�
NO.�p��g��`b�X��3͗l7�˺k^K޶iJ��j{-h�	G�(4O�ٚ`��:��].[J�%�����i@!��B�Rj0����y�������%u�߼/@1#2�p+��?��kD�B���<��(��O�j�c����WE�]�����G|��2�|F�ibD��L(��w@.wV^ŀ;Ai@�}ߗSR�s��a�r�8%ƈ�f�=Bt�)<B�ʡ� ZNnp����NgA��N�z��&�$��L�k�7>G �B<\�D�1�E�W)\�}M� o	u6����O�sH���c�1�?L҃G�b��e;M����<�B�������Z�m�u�|r�!9}A�.u�j�����}�Tk�!W��5����Z�r��ʒsGl]yhI���j�
q2�t�
(yޅz2v>��S�NA�c��J8��?b����
��œ �q@�ډD�VO��	��a2<��\*?G����K�A�h�ؖ[�;pǖ�1��i��$�MY�=��m_�q<I��o���,������˴�n�B[o��4�/�����O�T��^���ֹI�Q	�d�|��-! �Y+ ��s�6).V"�(z��

k�C+��
��K�i-���7K�m󋬯�imگ��j~F��o�y��F+)�?���N{FN��~O��X���(V.r5B�Ӑ��bD��^���9�q�r�VMs=��!��ğ�^�M?;_�]KHd �ї�i���:�3�?��)O"8��=� ��(�����<H!��ͳ1��d�&�<�x�]#y��{���D�BѼ^2P�6Ї{LaI�MH�,�Y/Z�ttY-�(��u�<[}m	�K��c��r[�(ɯ^��X
G#iK�gpX���T.Zj��6- ���6��zX�Z-���8�r�|������OF �����&�WO�s����3!dPuZI@B��s9��EPrՃ%�~�9����0��\�2B�:L�`�&��;�J�F,�t�R���3Ɓ/K�f�:Q5ʓ�JO�5������xbX����	cM��'��<�p&�	�s�ҁ���lY�<'`	�K<MZ����B��$�&��(6�t�kߙ�V�إ`�㼵:W�l�KƲ��&��RҊ�7��w�w+K�[u���P��!(|@yLpṄ��>i�kdS�k��Q��/�},x�qv����
���e�����5����	�N�]]�Z��U�V�A�H$72��R����x>N�xsf�K�$-�Y3I�e!�sK�#�Z��b��'��6Q��5%���+i���!e�L�������|�y[
ֹr]^���՚�� �,d���e��kť�h�4?z�Z����3U�������M��Z���y�۩z���/���@p��1��\���C�W�s�w ]�BD��?bƌя��u_Ӂ2��C�22u �N,��ވ������n���fC��{qg���//m�4o �c�5N�H�'7���J��\�� �i��:��;��
�.�����O?����BǪ�D� ����M_^�m���HT+�V疽��`�l�4Z��6�g�K���5r[S�zö��i�U7��B���T(-Pc)�����n�-޴ _kW�\���B�xC<�����O)!#!�y�h��_CË��['�P���m 7�K����������w�9 FP_w�sF9k+J�~I��݌h^���wT�,�<_D<�C=�\Oƕ͂�#����&����V
K�Z�ݚ`��[<Zﶞ�������֍Y1����k�LR��$t�0�1\,[�,�BoV:����wͧV0ke�v�u���� DKZ��J���Ρ|y������!l	 f�N7�e9-�������R䲮,ֳ �p)9����rz�FH�Z
�MٳD�8p��� W;��Z��Ѕ���rx�m��ȩ����
�Y����0��x_��k�,��i��*4����)M.�Ts<��^B�g�&9 ��]�,��5Dvɤ�.�HgMF����t��;r@J�,�T�D��]�'<��|�u���jw�1Z	���%��P��n'���é"�����s�Ϛ�*�4�yZ^jq;[J�:;!y�t���ʯ����:_PX�e��9dR�l��>Ĉ �@��0��tWï#`�����2��߮��@�j"*�aLcqhqK���J�|~�w�˯L�v�?�F�>����k�j#�}����cW���C�"\`D�w@�{c��0���]��1"at�:��c1�rW�He����)��G�	ѽ@����[�q11夔�K�dKa���	�#ZJH-�u�
eE���6�z~�I��g�����s�n�e�8�� ��%�״%���;D7���{�=5-��j�h�x�I�RG�8��#LA�Xi��u�{2n�Ν�9��~E�Sb����8��-��/.+�7Zi��g��/Ӳ�m�H���u��G����>��d��x���b�J���sZ!���8r����T/��{��0�+��Wx��8dlh�qL��-bw�!?C羁�p�!�2(""퐳CN�鐽� ?$�w����w؄�pD��C���;7��O��'�z#�;��ˁՊ�'R�sG �2}=�B��f����><����t���E1�פ�e^�T~�ϭ dY�g����ПeV�-�,���ΕtB���I�nkQ?�JS׍��ӊN#d]_)�[���B�Q�s���(w�s�_/CR�~���)U���sk����έ$��Z���r�l�S]]��9����V "Z��!�Ka0�'��N�v�X�|�8v�WT�sy]�څ~�F�"��qr]���RBv(NO�<<@ �F����B��Ϙv��(�(y�-'n:& �
��5�b����RT�sNxk��e+�K}�����4a�\=X�H+��f�����:�V{���2-��d��k�c�bZ}�ɪ���\����w%?2-�+��b5gԿ��j�5��'ͫ���۪��VөIS�Wȓ��E�С��$DA9����D@�� ߁�A��:�"�� ���'~S���u[�Q�^�"����o�{gG�#��Mˋ{>�Mm �8x��{�1��hFWP���J�a�7"�k�I�������:�w�~w-�]"�e~z	�̹I�z~�����=[K��Z��Ǳ�dH3 �+��6�/�mZ�tI��d�9��-���Yu�|�<,�yNi�_i�i���[f+�����5�ʻ��]g�j�w?��`sV9I�k6�t|�z-�hK�ꘒK$�T}��X�J�U�k�WW71=rB  �����z*.�u��ƾ(M���Å�vI	�FxD��0��+gn�b����rYM�[�<����q3��m�F{疡-�F�Y��D?Gk����㭥�䀖�X�ƫ%���.G'�n�����s�E�����3�uY�q�i�ϗ
ʅ�J��O:)�y�����ѫ����eȕ���ZyX�]������`�8�2:x�u� �4{�x��!�D�CĮDҤ=�"m��&_1�@H��: � <r|E��X,� � �bO)�W��_���u]7-��a(����;��n����x{�ꜛN���/O�ʁ��tZ>�r0���5!�Z	X�e�&K�Ⱥ��k|[<ʥ���$��H�ѐ�Ԥh	��QN�O�.(�
0N�7�鶴���Q*��kn�:�sHuM@�SX��j=���[*ٶkm ����:�2��L���w���\��Q� X��xO���yq9���?��$����=98"��H���� x 6W5�P�e���??>�9B򄐨�L�wIf�2��}:5�c��!7]z��  �J�"�)�M�^�ZK?����[���9�s����|��:�5Q.&HO�-��`��|&��F���tXu֊��<�$������jK�������Z�\Sr�
�%�,�#� ��&٧2?�k�&��X��V;�a�[�n��e���:���.&�3 �<<({��A. ��f�#���2���Q]�(��p7�ۂ\� GU��>t �=�;�ոb�nc����JD%��ရ�t y��
�x���ȩ^@@�h���Χh�2k��/Q\��c>�Z�� \ݠ��7X-��������%\$��Z������S�V~��$dK�ɶ�m�6�[|�<[�X+^yH�?K�K��-���2�vA��c�f	�)�xڷ�W�sm���]��b	�V�X_�_�tZm�W���%�����u�������1�M�q�G�T��W������y�?�2Ʊ��x���%O�6-�{���;���?��� ���^����r@k@�}���a����'p�l0� �#Ƃ�7[�9�u�N��~�'���s	��#�b7�)݈���4`LG���EcJs�D�֦�sn�ܑ�Y��fw���������ˑ����������i]�����@�=��%7��{����f!��w"��,�˔�R���7��s�q�����"$���i��]9/�˽��/��kw���W��\ǡ������m��~����<b�RT��-�"���\��z�i�E���
VI^���tr��nҒ��I
kɃVh�����j�.t=���n7��DT.c����+9�#�MF=(�»��l�wǻ@���V{�G��Ƚ�a�#v���u��#p�{�6�}��8d��0�����ބ��/�G�m�n�BJ�f����Q���mWC�.�eCV�yP؃��Q�it]��v�σ��`��/y(��,4���2M^ͿU^Qk$n��B/<�D+?~߹r���MOb=	�!���wn��$��ZU���&���=F�;1F$Z^���@�IXh~��q�A��G�%S�A��?[�O�?W?��ʯ5gt>Vy���fWV!��^�������iV�����7\(q��=#����n�7�{;1�#�ۛW~O�돽�ݦ?�~ȄGn�����6W��D���~�@�J0 �+����oW�s.1���ON��q��Ҳck�< ƅ�5�������wmhҖ ���,kM.kR�߬�$iw̵	+Q�ޖp�l�e�~����!ӵ�t!@T�R)�ЮN+WU�l��D���R��ǆ�}ݶ����U�Uk�殖��TIY��:o�A�O�����������-�xz{�:����8�z�;�FdD�� � �v@� x�臀4d��=�^J�~�á�`B,(��/�n-z��/��?9��ѣG �����i��� \��\]���v<���Đ�Yޤ%����t�N�o	]Kps>�\�/�OW'X(�g��W�'=�e:K Z¹EV��|�yK�MQ��l��_��Zm�B��N��-!��Y
N-�-;�����p����l�2m��\�.:��m����_�ųUf�,e��o-/��\�W>��),e��M'��H	�ϟ�x<���zj�a�q8��f3�_��x���qww��Goᦿ*v�cwu`<���\�}f�{l��
�m��WȀ�ƾ����1�k���	��U�\�&�Oe�ƥz
��e�ֵ��$����.A1-��"�����|H��FL廍��6�Ϧ��3Y�9�,��4��un�[y���I:a����:hEj��b{�|����cH��d[�V�j���]b���x���U_��tzk��]�����:^2��
�Jl��y�f�s��(4�Ŗz�m�H� 2B8 ĺ����~��;`��� �	�����4��u>|����U����~�!�?~��:�p���9��wwϑ�{l<nj|v�`V=QM��u����lB��=I�p�{ku����y\��F������?y����a�|	�x�|���Y���b�lk<�V�S!z�jA�y��.�^��
A����?��V���;�#���U�զ��-@��N�g��X�hN��N#�\Mx_�%�y�f"�=��U�/v<~�������ɩb��`8��c������^�ވ���������3��ޢ�;�r ���8 t�>��{��5<F�1&B& �D�P\��@��\�Zއr<�	�[�B�L<I4��P����L`>$�	��M�mM���%:Eg�sK�9�&�*����*��[��R���r��J���Њ�jk	�~`>��g���d�L":1/��"�ETSY/,Ƚ)���c�6��_ڴ�MN2�ߺ���8y�^�J[?o������u�O�8B�4!�G_�~!H)��<@7 l�bFp9@>���6�b���A��ؽ�% 9d��d> > /�{���I���sBJ�3�N�|<}��z�n��q��;p�d�{�a@���밹��rm�FD��)w��\Tdœ��͝c,�w7��	��-��y��~G
t疛�-{��W�o��Z+��j!_-$,��2dM4���iZ�X�~	��Կ�P��S��%�d?j�p~�B^�g�6�q�1��t���ڥ�jg͛�������'�[~f���o�]����7M�شƏ&]��O���v�,}0Y���*���x�wl6����w#���{��p�@x�y�q<���'���v��7�U��w�������~���������?�C\}��c8��!G4 �G����s���G�n���|9�K.a?p�NE��͏�e48�hD�w���	�_#�1�\FlWє38�'r	��Pv���,�h��s��Qk�}	��ϲ8ꪽ�U��.� �z� ��W��Q�鲎��z�(�P��4�Q��p5V7���[�1�)�H�P��s�BH���R)���t�� X��0��恜�Ih犭<�WQn��sJ�Y%v§<��$�b(b�����#�
5����Hi>K��\]]�ș�'CHiD"RK���j�Ҕ>w�g�ue�8�4�vaAC�PyK�T�G	��K����┑�ن��X6��+�p�~�S;�te�:	��_���w���<nk��q�}q;D�
�
n�+L ��S*ם��N�X�vuT���Tb��CJ��G�B9��G@ᕅyN����B1�!��pX�2��R<v��[� D;���;����d��{ ��v�0:��o�i�.<@B�bw��8���A�#@ϰ?~�}z���nv0�]`����_�n��������ݿ����(����>���o]?@��V����k�www���o|����ַ��w�ݯ����m��;`{ܾ �� ��F�|�T�]c��<�ٷ�e�&D���g�p5�[�uT�"��5r��W&qiTH��iL ��'�e�h!Bɋ< &����n!\]�o���*G��V��V����O��$^%z����H�W�0�,#߳���HޭU����P����H��E��t�s"�V�7�=޹y�wb�Ei��n�u�o�� ��~V_��V@�}�ct� ]���v��-�H'u(>��{�v@���aq)�0��{�ww!��w߅s��]���7o���>���)�O>�{ｇw�~���ٟ�͋����
�� ߫��.�o���_~��-W�����߸�o�Ɨ�{�K���qw����q �߇�ρ�1�������G�:P�1�[��Ϻq{�|�1�ֻr=��������.r���/0��7��?t�ǐ�Zy�nB�B�5H��S*"�s����r�� Gp."�	�P�M�9I�Y8����3U�\(�TY^�ut�>"���w%mF��fR6o�˃+1�3�r�Ee/'Į ,,�k��Cv�|�D�DD�\P/�2I�[*F��-'�6�([�w�� �	y8_M(�qP��q
!0�Ywx���8��<�tj�!P� �,�H(�Iх�6A��Y���r� �4s�wP" TS�X=҂��b7OF7��3��(\�r���>��H���c�\�!��W7u�UVw%��P8�O��rݗ�`�9q�y��ٶ\�����<���:3�����i
�G����Pn�K�y�p������]Y'�9ct{8�E￈q����4>��'\�-�n�|�bx���[x��p����c�u��{\?�c�����=~��~�������{|�+���H���xU�B+_��{����<���~��|�;x��	�|��4�s��q����х@:�xw�}:?��c�7���ߢ�MY[?��#t��ܔ;y����pss��~y�!�\���=b�����b�*T�'��p����D�&���в6H����,��L�Z4*^���nj7����3O�-��/�t4��S���3�B�0���'�]s��l6�(�r���0��`//F�1���k�u�{�`7��T����C��!�0�Y��Q٦z?H���a����/�;��tm6��U���/߱V��y?@���<�y����u���\Qr��e[1�9����fJi������y�sF���n��5�c�X�e?d����z���!�@��)���C�����p|�O�}�����6���}��?�G�3/~��K���w���f�#n�������C|����O>Ə�p���o���SlwW�O����a��?�!��bW&t&7:�a��x�Џ 
�b���T3C�t���f{ꮑ�,�}�� ��""��C&$�j�-���"�gLŶ�D�`����Dmt��/;��p�pH� �P��fa��깶2H�[�L��I�'E�D��* ����������e�D%m~�P! �p�"��c^
$�=�q���vc��G֏yq.!g��(�d�#��$x �pF�U��T�3a��W���]ժ����=�>�F Rm��P9��Q�@��+8_�7�*���uHu����
�u�䲟@5�ԕ�c���c5��Ԟ��R���S�H�%�	1�ƥ�D#RN ����W����@��0�=-�����0�����r� r�PõSQ�}5��!d��T����poq\7`�޳��h�qs�π���.���#��g��}��Cl7�8�>���w�ݻ�_��'��~�;����?��������/�ޟ�o��[x�Ȼ��U�k��8���
�~���ݿ���;��?�!~��?�'O��������~<b��'��F��=6ۈ�pG��v����+(e�pu����"��-b���Ï�!,��-^;�6�������NO�z�6G`9�[����z�٬�"x�In�7�P��}2xfAf�5��əY?k��2����O�r�F�9��_�//�����J�qˋ���{��什�Jc�8O~<Nl��Pe%s8�v��0���x�ߵ�&�s�K�ruz��n
�~�W��8.l�r�v8V��>�+I^��{rU�s�0�}��f�oV�.�z�I�+Ǧ��8�+ ���
��qZ�-���ҳ��Q4������c�������Op������5>��noo����O��߃�#v7�0������8����'������2qݡ'�~��_������C��[�����Ç��o��?qj&���څ����3n���������zį��|�o��x�����"�������>���p��ǌ�R��I�!cȟ���}��@�_�����C�<n0l��(��+Kr���9D����?�:]_­7S�f_�W��b����g%��d�ROL��'�^�Ky��'�,G� ,�Mz�`	~���}f��&���湨?a!d�±6}e�c��5�ςR
{ir�v#"d�����0Z��va�$��H>��NG1�m$����v��JY��n_� �P�qt����0L&���:@4�y5�l�[\UE���K��++����O���i8�I����#����2ƈ|U����5�{?"� ��p)��AÈ'O?����s�g�6���E~�!�>|�4n��8� x1�,�l�9$|t�������x�������F���?���~��'�K_���c��px��>쀫�Sٟ�ވ���p�v����o~��.����8���[��u����0��|�����/��*b��)�� ��������툻�;�𸽽E~ї	DO�<��j�C�T�s�K\�.��G������<)�y7^�ft�?,��-X�N9Q� [�Ri[�9�ϟ� �2�d�h���	d	\�?֨�
�|���n�W
����|n�?6�v��T�m�B?�\/�9�x�t\)T[�/u��6�+.K�J��6u����$�Ԭ�x_@���J��,���l7F�R���{�,�����i�  ��]�!��?,�k�ٔ��b���E{��r������٫E�׉�u��#nooq<B�f���)i�  }G �� �	94�����1�x�!���M�a0�����n�M�b	}�cw��W���Ę���.����=!���>���s�&��7�	 ��׾��ѻHOkT�WHoD�c�a?� �~g@�\�o�?���-��� ��}�0G�=�f1v@��p���!n�}���!�!g��Ce���c�����;\]=�a?�we����a���[xB?h.e�&�D�LڅM]9q5�-�e���z�A#K�P��VP/��z_�ѧ�(�kDD�t��d>�y����2/�=:�P��|�l�	B��K����#�ߚ>롞�B��]�-��VZ��ógO��p���2e�4��D�����0�$G̠A�H�s�"u�L��п�G��"6�ʹ*xz{�gO����6�<{��~�t�]��'�縺�}|��]�����z���`�l�1���y���p��q����O��8~������;���o��~"!�~8H>����o,C�������;\�n�ew���v��}�kH�����:�}�6�p�ӧ��1��t���C���C�:�>���d9-���ŋ��]
EI���E�(5���|��B��v���ӭ�{�*��L����K�4-��g��k�|���kB����ڌ�F�$�T2��s�;W����(�s���,���	�t���p{{;�E 0Ws����gK^2����?����]��g���?���Ǿ�<{����{�ۻ�������s�\�V�6EP�x�9y$d<{���9b���#|��_ů}x���~�����O���o������x�h������7z�uq���JO��?K>��8���W��M�1��U]�U��8�X�*!"u8�G�CBN@� SP?dx�A?�ͥp(��9ydtH ��;�����߇��o�7/՞����]�9��6D�N��{ zю���ߝs}� �ޏ ���{����{��{�L���⟦�O����=��/p� ���
�%�a��p��x��|"�{<��C8G��;���[����#|������+��Ï��?���}��g�s�!	��%���o"ƈ���_�2��څ���!z���wt���/^��������pw��ς(�4L���.���w��1�C�_7e\_�u	�~�1U���0t�q �6r��������W��W�@����G�>������H�~qؿ�G�|�������w��� 2��1r���?��O����obx�}�G܍��p8�+?V�T������������c�&~��t;�G��<yxk���6�y����һ����P�4��w
İܮ��	��1�`L[9�_et�W86�������=��=�Q���O�GO~_y������)��~����1~����/��/�ގ�����B��?�g>?B ����L�|�OO>�>~�1=~���d_������X"b�X}���1�� ��S�}_N�v�%�����r��$zR�?]���k�v����x�����w/�����[��⟠������|	} 8|��ы��!>~��l6��?�� |�����Fl��#����=Y����c�� �v���x,���;�p��zp�68e��@��p��c�v;�������{�O�tO?R�Ƅ> |�w���gx��w�x�-�џ����o�g�;���z�=�p	WW���+Ⱦ�ј�\__����6x��/l6�Ŀ?�ʾ�{��{��7,�/�����"����}x����~�w�+�h�������?vB������^�9�xO�tO�tO��{�O�tO��#D�B������G���=��=�ӏ��{��{��!���tO�tO?B��-
���1B    IEND�B`�PK
     ��/Zy����� �� /   images/cd711d72-4439-4fb4-bf4b-39cbaf4dbd75.png�PNG

   IHDR  }  �   �=:   gAMA  ���a   	pHYs  .#  .#x�?v  ��IDATx��i�e�u������y���G6��HQQK�my��Dq��XHA��P �Nbx@�G�	%��� �dŲeA�$J
%R"š�졪��7���3��o�}�{UM
QTmE��i>�{w8��k�[�v����q~������pq~����q~��9�A��8?Ώ���q����q~���s�??Ώg8���W�^��x��ſX��-�wt����`�>�d�������z�����Wt����q~�.��~�Ϯu��7g�9
d�?�A��ȃ�V����lF=P�]`'(����yI�(��o�usdY�2ufV�ñ:���w���]X^ �����;S(����m�s�??Ώ�G��q˓�j��R��i˳P�9kw��:@�{�xML��1��A���ն�x��׺�}	��C�1F�x��� �>|���F�4��E��%�́���*D�T?k��<*������w.k���_�k���o8��^����e�j��G���7o�H���<�:��U���!����������9�����Q��n5�����G�-~�)+=ߨ"��&��'_E�X��q4�µ��1:�~�$�������.Z�-�}���r�me�E�����}"�Z�9�jº�T@��Ԋ�D3�%�0�O�wj�q���Ҝw6_�'wy~���E���"4�
ބE�/��6���:N����dǍ��ߢұ��*��¿}n��>?�A��8?�͑=�	���X��w�����lB��S)�
V�c��K��8���9������
�]D��*��E��kp6����|�S������˘Ň���������\;��Y���NNE!7B�#�`Yoc�����T�w-c�ۼ��8�@��Ǩ<�\�]B�����T�XjQ8T4��@g�qce�Ca0�w�2^�*�<�Ba�|g�n�x�qԚ(�-��ʵm;wv��h���8����x���܏�~��/����0�1WW����B�_��K`+ɞ��?�M�m�)�Jw{=���i�0t��o4.�<�ĭ����)-�
����N�\�V��Ң�5���(�˿�}!�u���<��qw����O�dVO(}��\�����<0����HF�R�P5����{&Vϧ��QRAŴz�b��%j9��q�Sʵ�B)���*��C����zh�7qr����������3����?^9�]4��5!��'e�����~��IJ���++����P�G�����eWQT&�6Za-�AUH1[������h��w�Bee	ɍ�d���Gmu�K��Мzķ~��'�9'�~u==��+���y��X�'�Aʐ�[pʖq��#$a�5��_��uB��Q��Cq��[��c�V~ ��h�/(0��
��0�2��f�<V����"Lo J�R}dy�������LA��:��������n�WYK�P+�ie�� ~Z�o׌�Vvm,�~��G\F⧊i�<�=���� ���]�<�lA�w*'���Έ��a$GQ�/
�a���:w��vM��� �(�̉�E!���C|����͟�_���
�P�M���sC�o�x��^��m��XI���������dw*g�@^y����}y�����_�����|���YT��2)��@V��%y������ĭ�W�%��e4Q�e6�S�W:G|�
JaI�P�.i�
�yJ�ja���Z������c!��z��D}t��h���^m���W%O.�7�����Ķ�5R��{�L>�%?�M׊Bd�i�{4>Q��1#4Kv�a��N(��P�.�m*�n�C�'�b���էY|�O���'�U3?Z�O�+��8�������|���f�x��g�PPN*�p#n�#Dd�؁#��E�@��\֮����_"���l�~�"�5(�a@��D�ف}�E~t����穀>�XBrjQ$�AY3�^G����'A�0���垞�T�n���' g���]���r�ړg����'����3����|���O��sByV��5&��w�"��QU�~���Y��=���=�|Зu*ߕЇXE{{{�f�:�
^�|�Vy-%�����>�Xf�D�����cZ��K�ޯ��/��Z��W?z���'?�s%��R���) 1��ʆ�:��3X=�Px/��a�C���~&�o8c�GŁ)��i�*�ɒ��,�jvG�!��@�a!M�sګ�k�1�Zn��� ])�%�t'�k�$*n �ؔL��A�QЄp��đ��#s��$�:�'n:ً8B#��4�	}tp�f��*��$	YŗO��13�pj@LR�򥏳f
�]�j�H�Y��RQ	U*�"��YM9���6�U
T~�E13�T޻C;ҨܠI�K�׆xo��2�
)�!���ڕ2�C�׼ x�8n~���y&�os���~z���b�����������2�-l��ao�R.�b>�r� fQ�vE�U��麨q8���w�0�e��W��	�r�6�9'9�� ?��6-K�� 9�� h圌vlHF���.Y0�w��#�7(Ӕ�d7o�>��d;��w�=��I�<��+>+�XJ^�bq����+��2𪵂-�$���Aq�0ĭU	�:�����`N��"��5Y��5QŒD�%P�fmU���)��,%�I�pm��C�؀���CB}���ך�-ψ%��jI�jB��*I�
�y��4v`g$����5�^pL��<��0����I�=�6���C?��j��)�Z��=g�!�!�T�dv�p���F����G~߀�33}9*N\.�X�lƤ�(��!ͽ,Q_�S���ܤ4�a�z��GFD�TKe�b�m+uY�r�Q��4�'4���H����,�l�Y���1n��t)zo�;��z���X�,^~�D؉�T��Uп�V����-M�+��9-�y<�h���`{�ʩ2����vd�Qpm���sbJ��M}VqkM8s���2��T�����:_�>��"��Rh������P�^�/�p���U.�>�=?],~,�8�9@Je�Zx�p���}��L�wS,J���$��5=Nh�d�m㺱���\kqʈ+���@5G�9	���4K��9���W��K�6�h��(�ʜK�p�œ<��*�t�b��>��"{����L�G� ��p��؝���=���UN$���W�>�*Ͼo�OJ ��Q\�����`ǭ�~��s�E��2�Kb�n���g#��=�K�'�MV�uc!�*�Q�$�s���Mf��9b�7���zM�M+���HP����&.��&�V1	ٜ��R2x�}�����݀`/�������
񚴾B��C
mK��g�}�a�-=���d��T>�����(��e�^���O�'�-f�~���~���X���6KC3��PR��
�6�_=�A��~�Rc��Vq,j�\�eS���A6��7! �ϊ`-��p�Ǖ�\��dsAW�'
�Jx�؅�{�����J�gi*P��࿹/���s�ɂ�0.���fa��)3a�Y�hPO�,�[2�
�� nC&������h4y��n+�h>�O�'D�q�|�����^(V�yO�����F唓	q�gd���!�o��;|Ow����
���F��ŝ%��C�W^_��&#Yۤ�н�+XѶO��k!�{���I�^�į��e4�����?���2����?���w����K��k{y��⃟�h�O�L�j����$Ǉ�s���P����w�Ȇ�jg�O���M��F��k6WR�.�	s2w��Xd��\����%�&��!B��DQp@#~�[��c8���� <�M�?�p�3��5�[G\�$>�c��";�����y�8F�ـOKd�X k�,q�sw	��~H���O8^�S�z��?�Znm�5]�o�����ִM�Z���R#������{�,��ĵS���-\M/rycR�`QʷZ@��%JOH��j���]Za�$l{b@�c�PaT�6bZ #��y!
�X�l�Q�b�	��wl%�_Ę�B��x�n@����*%��r�WPLeQ&{�.�}DC*�.�؃_Q.8���-4�7Q�N��W��_�x$�c���54
W����߮�+��u�6�W3�΂��"0�q4ƌ@�e�LSZ��`?�L'�fa�� ���vs��47�R�-
�|�*c�ɜx�[���\Ka^��Z��4�D��U^�i"v�]4&�H���՞|��ko$$@��kMy��R1�L����ָ������b<Vᶬ�SL_�O���UT��iPy��B�̆J�<?���T--��6��3�]p\���K%ZV�n	�Tf?�d�Vuz��S���k��K ή��V�-�/�@�f��=�j�N糭�����~[��"O�ybu��?o����-��dzhM|�;�{��`|x��x�~2�o8n�7��#�9�C�:�A"S�(�T�f<�a:��.ǡRks>��ϝk�N��kL�x��p�%�������X��3�B�+#��?�YB(�"&ez��ck���\��c�)��kamm�����o���0�ֵ�S�l�E��k��0��d�_'�����b6�t=��d�)*���n���j2H�29�'�2�L�<X��)��0��>V	�6��tTvu����.-��Q�Z�)���%KRfo�%�i�\�����:�e�k@d:o�e���L��@=����G�S�EL�B$�,%�a�L����,�����P/�_�('�&!�[,e�<��N`�0����=��6�g
�B`�e���V��͸���ԵD�_9�VI&ZT>�<^oqp o�cU�l���#=� ������\)<��'w9�c2�!�nhX��'u�w�F@�f�h��l�A�������I��y&�\��A k*Q_`���u.�8�	5��=T�а=��$hr�[yM{��!�����}�J�@�]�֭�5�'��BP��^p��1���d�DxqI=��P���ҋa���t�21X>�� W�;�����͙����h��{fu���$�B�� R#�Q�i�2��^��NF�1��75L1E[�b��Sf?7��ȏiQ�ix�F{V��|�_��6<�0S�TH|Z���t���M.��4��~��ےF稵�f�;SAL�}] 7���p�B�U�ֱ���l�O��[Z'�{.2Ւ4.��t^3g�`�j����h)VZ؄��*�3��� ���W�x�f���j���v�!:���V��m�����X��x혓q<WC���:��^��x�'+Ѡ(=��_��Ƿ�󋇑ϜOP��&#(�HjKK�g��L�<M�ʧ��+���rI< @zUt�Cz���&u�n3\��E��zT2�4�l8��>��n2�Q�l�v'��Ԁ��%�Ŷ������sy������SY<��x"�����)鑀	��Z��$��S��1�2n����q��Id�=Ew7,�n[�vE��Tc�VCl&*Ȉs�G�v��3��5׿]iWܮ$ ��ҏ'T��Ǵt�9�ͷ=~yCđ
 
��R��HǊ ��g�*�uz4��uG��*��9GB|�H���¢8���`��m>�+���Z�z�b1�!^XiMwmZ���{GW�A�A���g�01�Q<h�������H��Y��:'q,
��?��ĂN�-�"�I�W
�jK*8
�ꙕ�3�~ƛp31��u	d���;NS�R��y~��j�/yȲ�R2e-�6���&���͆��1�78M����F�s�,��򚰉'l4��[@�!��Ţ�� *�q��5�����:�e2�T�i�%��T<��� �hP	�ʦ��2I5�i?���긘�G>��-^���H�:9����yI��ڪ���S�ejo	��g&s�et�(A�-|^�Dť������-��A�Fi��ԙ�8�|D��v��	2W���C�#���!x����p$�� ��3�WQ�_ai2^�PjfX�$��t�9��v� h7i]p,i^$���,<ǜ�rLc'ֹ+�v8�v��0!�M��|��c�s&���]��V�@�������
�EΑ�p��D*y��7IE�E�.>x����	�T��J/P�8'5p�.�!����!��į,uuؖ�/}�X�F&P5
<lnn���Ǡq�{�0����/r!�d��Ȑ��6յg���$�l~�W_[OO�5���'�r�|�O�a*�f\�����u�ܩ��m~�9�s�j��Ϝ�7޿d���d��R�)���K�o*����j�g��A�f��s;1���/4�q4�sm�9^.z��ʳ���Ĺ��)����3I�Y�$�[�R�U�E��][<�UO��D��r��E�fj-V�����\�f��eM��ڷMMDՖ���#'�OB
���@�+�-!�Z@T��ǵ2���"�%�)n##|��t:�\G��;��zz_�wu<��"�C6M5�I��jہ��T�'bz ��8#�gS�.�畵�p�k*���@		�*As��>�(���uc� \5ĉT�`iJ[h�-���� �� ��"�=ه
*�?�/occ�o�y�7���Q?R* '^�-�ɻ� Sq���	5G V�_ ��T+$c��!�B8�!��>�}�)�R�h��z�7��nh,��h-���^G}����I69E�Y��ɏ����x������@t��i�ke��d0�c	�p|�q�R��>���Oܦ�U1��%'B��I��I\�
{Z R��zwkƹ�m�T���K���X8
Θ�^MUES��8lS>Vũ��;q`���d�s�窤Z�!���1�����s��i]y�21�����T��ѝ��1Wzc���m��q���e*	��$�(@РeUDT ^3�pɝp�@�,��&�Q֨ʅ(.�$�h��v���
��s�K}9J�����V���Xj���f�w�J�J{B9e�vR��%iA�̎a�&�R_�q��@%^r���=�>�ZU�9O�|]le?��Xf��O�k��W����d�9c�\�J���k!u�cȆ|Pb]�F�PZ)r�ƚ��[��]�&$��"ZޜD;�q@�5KZ�VF��iu������ї��ck��k���:�m��9B�Z��A�*q3�^\u��x�����ڞ	����D���#�A�=S'0�b�z+��Ͽx�VL��x��7;�@-����q���ʢ�
~�Ų�0n���|@��6?'7��XwH�H4���>�=��R��C5@�IB���3�o�ǳ1}D��FTc��Ť0QaP]+5��d�0Ƞ�d�کf��@��e�g4y�)G�,Mο�8K����q���Tz͌���1�!���Kj��k���ti�^�=V�3�F��Fn;�Ť�j�Z��)Qߣ\�����XRP�F���)��5ݠ����i�l�d�\�Uf��¨g|6�<.�x�M��8�o�x���S��X�
gT���rC8�	e�ATa���7�:~@3Z|��ԺYd+Z?��g��zf!?VƌR��`^gk�w]q��u1'���y�Ȏ���E�������d�b-YQ�Y���J� !�~�(U�W+f^g���Z\��Q4��Y��X[0��B�2lm���Vk愸S,�Y�(����B���7�h5%#,���V�Uf+��tAW�mRS��;s1�y�J�"�����zIf���"C�]E�R���ٶ�k�S�ƪ��4��4�.r�:�a"wK߻XS�NT���'4׉ u�(4�x��o�K�`�����]b	BS�ک��v�Яc����:&�֙L�m@ߩ�U�q)׵�)�X�s�e��ڣUʛ�sN�\\^�5y�S�2�ڵ��g�}&v���-����J�l�,�hY|�p�t�)q�5�N��J-�5q�$��<��Oi�pԊ��"�QlbE_��#�V�8��x�����K��5�%��R���c* u����P�i�ȸ��Mm��%�6y�e,��LT�h��L�
��x��@?"�����xuU��qs�yS�&�P[!�9d�~�G���	�(�ymO8��% �u���&4��<��;�v$MJ*�B�K�����*����������{D)Nf~�W;m�vi���8��pr�n_�MN0_�Q�)�9������D�4�,G�,�t,�%�暠��3q1u�3t�������К!�.Yn2w� �ν&Ƌd�CF��BFL�5�s7O<<^]�F�O��h�Iw� �����Ɉ5/�4����D}4�&�xR�F�T���"���t�������+g����8*HbΊ�1o�r�p�Q�˱�d'.F|ޘc�Ϛ&0�M�\>����iC����B��4�cLA]�f�����o��x�o�A%~Zq�dypl⩇��I�8Ӗ�ዿ��gN67�2> ��c����#�R}ZMq��hM������h)���s���2&�zdwq��b\��$��JuXD+�����&T�M*�2�i`� ��T�z�I=T�2n�e��(��,�����^�k]�ޣD-q$d֑����3���뿝���,�J�C������g�֩~8+HZj]X���7A�u�ޜ_�č�ՊF�����%#m@�/11ߣ��-͹W���HAy��YI)�w<�b>���T�(/�&�"�9ܶ{�kd�~k��9��9�ϮA��5�5�(O��L1�������&vY~:nK���⪱��GT6\ϻb�y��T�=5�(�wԵ�nW�7o��	MG�Q�׈�z���X
��Bm��p}T�B��E6��c����7Ds�|�S���G�D5��>3ٍ��
�&>��@_W�LN���B���)&Jr�/��v�n��5���	��%��6��
j��q��@�T؉���2���,��d�<�%�g	�	��<y=����������ع|yo��54:��Ɔ�prc|2P�f;���-ӿ45"���S�5�b���>�s׬cee��G�6V	|�opOY�lƧL�����3�՟ۓJz��r��� ��Xi�{��K��7$�N��x���a,^��j͛�����ss&̚cV�}�9���x1��Ek��n�s��Kpk�6D���Y�䊅�aQcDH�ڤ�J�������D�4I*}��?��&�79���|rS����I��H��|�XqQ:�m�B/��43��dK5Z�7��ru3���8�%��b����EW����ix��lS@d��O������tO�ȢN��gQ�ҫc-dqE"H�"��dH��I�L����!�':�-�2؄��P!.a�Ym���dq����qV)���/�O�oa�-��A}��|����S?w�$�:�!�ȶd��JH�}4�_}˹d��Κ��>"�'�4i�FpAB:����e���n� ?{�Q�N�S�H$�9h�����1�r���	��V��-�)�tQ�^�R��R'�aR��v^��\�p׈+��%��2��!|>X�d�ߧCŔ�3m�!�����=�$X��s� ٍ��eu��j����׳5������Nl
���.;�ws<��敪�ޣ��e�̸L����$���?hD�,���I��C���P6�0��d��g��D�i9�D��Om�[G�l�e�*o��M,��K.(38�hAؕn�s�5���)~�g\�|�����=R&�j\e��+cb7�MK-5o5�Nm9��F�B-����
�J��(���$3�	�A�}iI�J?��
�FW'/%Z�|;��,�Yx7���o��<����1�����	�r�Zh��П�*�f�x���	XS�E��e�m��α7�K���Br��]��0��Z���J��^��	X-GS�4��j=�~�G��� l�
� �*_ۘp�G�] �AvW���9�B��x*n�&���|:�'�S|�uZ��	�kv{��ʊ2��S��R��jl�2�I+���-�%�y�G7�M9�⫐�A!Z��L�J]�KÁ���T/M�z��P�/��Y��YuaP�E��u!��]{Y�S����-�-/������#Z�Y�)����M�_qʧ@����}�#��p�>@\M�y����O(
k��j�x�M÷�ն����y�4���4���V���T�X�=Z�j��+�uğEQh"DƵY�$�F����J��Ljk�㛖�ر�M~~�FX�_?-I-��"�i��r����[�LgBbRO枟���ե"r�u�,^k��:5�q�|���Pھ�Y�Hzĥ��\�dDKd.�9�����\ZqDh~/���|�E�R�Ƿ�����մ���|�c\v
&�2��\�%F�F"b�$�[�����>3W�A�8I��sݰ�.���x&Ч���"���f�GA��Ɣs�{���s�9�^?i�^I����":9)� ql��u#��̞��K���6ۮ�fv�9�P�\#�ʦ9�@�V�G��7*�J&�}��p����M2��I�%�������Yl���<5�w�w�u?^�%��MXg.-p2!X3�HRJ��a���/�}�����[z�I,�́��C�V/�£�$�ĺ��y�.]�	���{XݾH3��c������~�]mhWc<ZSA`�_}����]Of���q������00�Ǯ�
p������)s�xt�V��7����������,V�V%�8��vw}TAH��`f�&��Ͼ���W�
=�;��t�4��ˊ�%�T@�����)��v�m_�J��{.-�H�|Y�E�~�O~�
s�����9�Nz#�0<$�@h�8j�a��v )��\�GxJ`�j�%��������|\��d*��L���4	u�
1���*c�[̴g}�	<*�kkk8<��`(��lש���h�,CLjK�G�}q��~Z����1.�~ҧ]��M��G��@��kl����âf�~}�)���-,����J�|Iս�:Ա �ğ��B�$/�Re٢�mn�����qo�g �����n��ic�2\r�]IeM���]��bQ1&F��|�k<eb∮U�ɭ��d6ې����Z��gY]u��xw�����ᡒV�a�E���������2��$��U]QRA�=��YC�m�}�=�\�����CL2����cx�1�L<n�d��w�y�~�/_�#%{���S\�����k��L�dc�lvD����W`�&� ��H�hN&W�U���4�]]j�J�%c��]>�1�誚ڎddHV�,$�Dр˅�HMzS�����uj���+�)q��ro��~��U���`J�E�o7PL"5�[�K���Gd`�9:-��%�Gd�T�5��M�N�gk�x�J�"m�&>��j�b�%��۩L��T/W9MT��d8SSϦֿ�����[�Y���s"��.R��j���i����^��	z�?��o����|܈��s]�~�䠧�	�;�|��^kcs����{��n�K����V��J�W^��K�T���$���>F+a�޽{/��Zݫ����:��+�ޥ���A�F�f��Q4��:�K2vױq�%��'���ʵ���#��s�����C�0߷��_��;�9��O*�5�؋�9^�bl��|�
�#�ȗnR����GWiI���l��r4�"tgX�HqM�˻.4��N��%��F�p�����b��� �mؓ�N(V�/=R�����_��T&�Qi,����!N*�X�Z\�b��Z�'֡�>�v¹N�.�� �����'�Y�VS�˳��v�Ӏ/�D�x���/�K<u<�=9$s�M����$Gށ$N�5e}��!�v�m��r]gu�9�Q�ټnV�>?�J	~b�X�*!�:�!� ��lIƐ�x_�Q�$��&e5��4AJN+MHۑ��+k�i� Y���ފ���:���``��G���'��.��㻧�$��V�r>W"�ws������27�1*��&I���T��L��f���9�@��=IU�4{;%\�T�W�q�'n�t�)�|1����R�L�;�/Ӓ�>Z����ҥ���H��gb��(�TƸ�����s�d�^5�ۛf���KG�~��+�á��e�p�X5�R�M橺~�4#]����sj�T����ʘ�.�9�cR��z=ؔf�����B ��իWq��]�h�v�j�^��Z��h�ٗk���l��_�[hUn�� �GoJ�%CH�oUl��Y�1��ɧjUX�y�&���LG}�blm�	��pr,��mZ�\�@�K|�"ܭ���8:�P�5/��c��9�1BR��M ޸�qR��T�~��
��5`�O�x�8Fc�^�7�5��5��9^%�yg�/��;o�X_U7�A`��K��ƶ]�eE\���|pp���Kd�	B������� ?�ӿ����?�Ƿt.�9�SS�IC�"U�:[�Xkt��u�-L��|������cܙҤK��cu���\8Bkk��0��Y�"#|a�d_Mx^�n�d���&�4��4eT��\.�P���a25a�m��֖�qL�L��<O��?"�_�C�!Y���wvZ�Q�*9��׾կ�d���2�,�:{�z}�זM0�MJ瓱��ބ�����{�m-�J�ئ��C��-����:2V�2_֩�����*��Ҁ�5q?��S͖/� 0/�c]�P��\٥+?�)�te-�i�dq�_7�њ�ajM�Z�ffZ�;�֩��I'�3��l9<�������ʰT�Nr�u�jE��;wLK��l�~0k�&���������#e$d�i�R����N��]�0�����^�3Ǯ�Ӡ���K�QcΏ'�T��Ϙ7�ُg}�����@����J���1O,�H#
"�a6�C9?F�a&�-H�Q�b_;�I�h������yƇorѽ�W�c.�n	�-hj�Rd�PxE��w��mlx4��C��)^|�Ƈ?uG�!>�kf�;���Ʉ쨋�ё�i'J�(PI�@w��$H��(�$$G
>��Sa��Q�L0֎�I�0��+Z�#S�h��E !��@��*uaesI����:����Ե��eu;Ā�?X �,x^1�;����#�P
KZNU{�+�u"~?����lʄO�>��_�ݞ*��ɀc��G�\�Vz��"��}���}|��Z������&�/��?�7&����U6�����'/�Q ��o	���7��q�G�Ɋ�ON�ӷV�w<�f��1h�s�������}甆��/h:O(m���}u���Z:�<��у�b�ZD�c��������M|�G��ۏ�$~��E�qc�������g(Zk��u�W͒l�ˋT1Z$����{�eJj�llggnG
�h�u��Kơ�I36+.եQHlA���5�LlO����t�,��簒��J3@�ŌJ�S�Ȑh�O0��b9��_��m�^������Q���,����������4��b����ƺ����8'��_��#Q+�JL��r�ܟV�.S&����:`*�G)�Y����v)�Bz���v��t?
5&�Iߩj���ɑc��S�=j����i[k{4�B�h�8�V�.a���¸{hd���j뀋�Q!s���}�'!��1�^�&����R݁e���TLB�Vʞ>�3�G�Ꙃɝ~~������<��n�0��}���u��7M�����7��V6-�,�I��j\����&����'}|���siizݬ�eo3I��v~�~x�����!��4{B�
�jD���{�t�|��ױ����X[��G�/\�e��ߝ�GZ����
��W~e��w��^j��)h�u���I�4uݥ_�"(8&�Hy�l|�$�����������H4$?�H(�[i����:o^��(�kk\ �����芢��{}n�7�M�v�[�uSǨ�.j7@A����_�,�{S�R��s��|����H�W
M$�����������}�_�����������|η�\*���⍇'���aL��Z/2��<�X�h��r-����}��s��߅ďפg�g���&�+���ղ��Tx�Ŝ���_l��J�1:P_��R6V��s�.:YXY>��I�k�(y�b���ֺ�ݻw�/MO}�7�Ь��E��?$3+(+1Ɍ/�Ƨ�xI
��tR7�!BF��Ô�7�9�:;%�	�xa�����=��h��ۼ�eu6�4KK|�r,��O�n�>���4��Wx
��<��?�$�/�yC�+�P�c�ǌ�d�,�3��/i�	׸�r	�&�2�\Ga�B2�
�*��2�l_��l<�{�'Y�G1�1�kPb���s*P���4��b�th���Zl�N6c���5���5Sw$�3O4c��w�z˥2�A �5�9dM��n��x!{3�Fc�eT�s�������"7���J���,^��(C���|"���7+ur��k7��d.�h�o�?O��=��xf�w{W���AX�hR�tATJv��(�⑖`K��n(�޲2e��b�F�!'�Z�wN��R*����_ýw6��~Zj��BIdW-ɴI%��'{*��l���af�ԸU�1~��wq���\��O6n��74jfa�A��c%�͖i��:]L�s�R�Z褆�	&ajT���"�����e39Y��`$�Kz/�6���P(Ϭ�Nj������ӆ6�ܠ���0d��*T �$d������L�؈�`u�P���}1��}�gp啫��/~?�&�<$5&��h�S��Ϲ�m��\�Ɵ���ܹ��}���{�5���W�������D�$]Q��
t���m`�E��7�ko�?O����OC�z�M��	�t.�S4��v����C`�Ͻ|��?��G���gc��u.�Y��*u��fP�zYț�i����]bob^����%��}��18N��[�T�J�)���\��s��;m��b�繘^"�ږ��m�	�#�Ѯ�F(�nC����8��-'q;w�
�����x:�w����k�B�����:�8��E��o��2�1Y\4�^�1�cIF��x�ɤ��V�ˮ�V�'���<�:Z*��2��I�dK]+�i�k�T8	��Ⱥ�PV�r�bQ	#-M�
�1|��/��������6�n���k
���/o�|.���(J��M�rɂ� �/'�4��X��S���l�.c�D�)I�̻�3s��2����V�qM�f׳��S,��8��E\�%�,�Z�>��N�bPвw�>Ni�˦er�g��8T�v�t���cw����D�e�����9 ��4�=2����I캆���}k�K#��@Z;c����ƦɊ��|�'|U����g?��W^���?��J;Y�����Ģ�_��)�0��|�	��ߐYլ�Wg��g3��Γ��b��x�\��<��k�9���u��4h�����ܹ�g�~��o��h�5�@������i�|��OF�&p�8xa�Rt&���F�e����l�5`��L_�n$���if�vN�Th����`��kk=�E�!�#�斣�I�e1&���X�/��s��"��8ܗ�HO�=-�:�q.YTM�~�7^ǅ���+_���6�M�??������⟗�j�Al���w�� �Xw���x.�s�$ߟK��V��~�ו �fB���ߺ��h��d���:>��/��Np��w4�E�[�fo�4�ؘ�}��YGU���^�����}�w}�/t��������.�)�Od���ɲ���v���o���~��Ec_b*�s�W�nħ� ��$"d|�K1�9�|v笣�0J�֠5"��F␽�[�M]�0?�+hFX.>qS4����-<�ҫ:O߸Q�2R���3I����i�T��Yj�oc%��15�,-M�Yi�(��vKz]y&S�\���٭+��S���,T��T��l�<5ջ�֕}���T��f�a�~�ϻ��ŋ���nnjt�ji�q�G	�-����V��8���hFk=���:���줆��E��%�&m��MS�(ߗ5��H��H��H+��s�3��Q��>�'Ϥ�[�5��E 2��ѬßLL/�UZ���� ���%C�������} �hct˿�=Gl����ʹ	�c1yƣDM��\�ߓ���)�I=����	楏�*�NC��)'�"z���'�L(��l��J��b���R6R.�h�Z��o��ƅ5~_��7��� Z�X*�Nѕ����n���ÔF�JG*cŏ�R�"���
m��/_�ڪ���{��V_>:����nui����'��n�@�k�iS�Ӻ�SW[A (]�8$ßH���F������n"��Nd#
Qg�l���������8c�M'dKS
�xAŸ-J��s~��v��	�d��=^��f�q$���6�op���NA�8i��w�;A��������� [+��@0^`g��������#�U�����5%��\M�r����FmM��QK��������F8�:={M�h��#�JtO�=XX#dR�~��f7N��6$Mt��q����G�u���W0[q1�Ms�H7��M�����\B�^�?�&(v\Ddyr�>���2) ��4��~�+T-2x����k�(C���ca��QX���yWi!hQ�������'/��m	��*�y��(���F�.J�i_�(K���Ӷƕi� 
A3�`�y�P|w�Y�Z|?�;� 1�-ӗt֞�3;� F�
0M#��h-�pKW�Ta���ť�ї&wEݔ�6m,*c0��U��L�tzpkj�];�����E7�Z����z
J�!m�d�h���Jd�=q�H�]Z��T�L�\?4��hK,k+��2��h�b2�4�2o����N�2�WC	�sMHL��<�*p��ZL��!�Hu�4b����#��F�A�i	����X���ڐ�V�����I���#�@��uN����9��s���	�3�	�/�B�h�!���h7W��A���ڰK65�ݪh��6�8��_�*�2���UղR��j�M��_�L$�~���|Y2=�f����ѣG���A�9��ޥu�Xn�V�.pxhzy�b&����M��z��v�܇�S������&�=x��W�zK5���қ�����ux�r���(� .������lCX-�vK5��hgM�~K��$rO�����,j�
�aN�&|阘�<vf��HfO����T��<mV�{�&;BX�h4�w��`gs�2��Y��{���,��|3�2_���p-�W�j�j�����E%)�[[�}�H�,�&���la��䜳���8eI�i���#��@��-�We���H��\���T������m��%�%�H���ï��C��ｫ
@|����O�kg���-7L��a:3.�2Ev��vAY`�yd����H�GZ��qZ�-��w�T�T�r��c���k�QD"V`�g���/�3	���u��";c��b�N�9ĺ�{�]�HĲ���	��T�)0��6���p���g�!�Y,"��vh��JS3�V���K�lӈN2�䰤`��&��dg�\{ݔ$1e��e�Wn�������e-g�L�����L��8X�s�#VO<C��cS#d,i3�b�JF��k`��0�jp�@DVNn��@Iەq��,ٽ�a˪�J���]�ØN������X׋Tꊷ`X��2�qxxh�AUk&נ�.b	>iӫ�~6�Os����@@?	v�e�QX,�	��ž�Nv��Ny�4���M�]��0�-ě�����DN�;��A�t.m����O�+�l�o��s1/�q0:Dg��� �̠�+ݻ(*��} ������]�%��4����]̿�~�#$�VyK���DJ�eRQ���\$O2�_�Y��E�#���X�����2�T�E�Gα�� ^�m�f���l�.��t�s�L������z����q���T�H�>����@b�0�R�}D�~�О��0J\͖nI6N0������)��Mp�����l7���/��=�������6tSٜF��Ml):���[j@Zbs�g���#g>���ZwOwBZ� l���L��\T�*zs�&;s�٥DF��On6t}�?ƄE���o�[���_~44���wmL�D{�BD6���n߅�V_��X��`N�-���w&�h��t��{� 9�!��yG�]lP&����C�/����8_�V�����ޢ<:ڣ�I���n�y���������*�Vy��&���	E���>>��79�C��ʆO�&��Bʅ���f��@�ɩp~�4�
�[�ta
%���4��EN�޷���̀��rtújKP���ie�����)C��g�P�+}�Ivh^���G=����u�v7�/���vu�ד6�Z��#;�9&!�vm�U W���q��� �b��Ҡ��&�x�ŝ�_�*�ɣA+m��:1��R6�^��Ml�UVK�+��
���\�v�Vݺ�C�� .J_��y�T{w=�6�b�9-��� ٞ�Bl�r]�W
J��̻��h��aF9�݇��%k;8|�ר\.X3|�����C�k�-Ap��+Vo�Oe�
];�
���iNN�k���|��0�s.���� ����?��ſ�������D��.��J�,U�/W�X�٬8��F6�z��Ƈhz���a��0A��2]-e�ɦ<�?�(�E�$�8T���ΤI}��wz�y�B����(	I�$az�^KS��Dw:��4��m�ϭ���3���W���GZ�\��ܴ*�+e�ҟ�8���'����(���	�+�N��^Oذ�r�@�}Q��� �ZY�xs�= �^2�<6G�R�V6��OK|�u|�V������W~e7i�lnua��3P��J�(OJ0��+�ӽ`M�O���dܥ#���Z��n���Zy���������/��7�W9O�_���^��yٯ�k������Q�%�l���G�Q,=�6*��|���6.^��o��}����(���4�Ͽ��x���EP0mY�z3��,�$���7�_���3e��~n3��"ו�`��CZCEZGG��1�m%�C�27N���V�ڕ*?�58۴�8>��=������ ����~�f��i'I��9^�NS������������?���h��d�	����zIcӯ���u�k���{���|�
VC��vf���Y�rW�*�-�g��cs����D��v�K���k�_ǜ�#'���3,�Oc�*O�̥5F�wQ�O�{H3�+���1u/�$�uH�X�,�f�V�Kլ�~����8������\�D&�@;��g>���1�N����/���=gz�M&|�F�r��&�r�{�U�Vɛ6�R�,��p�}AŎ�|[K��>��@@_�894/�E�hs �z�hn�p���iД�Qs?���}6�,!M���2m�,�y0��n�)ˎ5d�&|
A�s���\E_�`��
p.V����!V�_�����VT`�O*�*��l��+<
s*]4�,��@hk`fNa��-�T)���kvכ��{r�jA��-���G�%����w��]�c�,�h�;Tִd��D+��Dӑ<*
�/������f�4mg]m��Ӳ�!8hn��#���EaL��)�(S��k���G���"���^�	�ڋ6�������K����>�� ��`+<BZ����f�ƕ��N�B��x�e�H��.�S����wdc2U�����1;v. ����J����O_�7�y6���Ct���m�C��"�yצ�`K��\��Ke�=]��K]�<₸;�%g���1���E��k�ο���e��>�U����@{������9��-���x�ZZ�o�����w|�⹫�g>bxt'2�d���B/3�I��h��A�����'m�A���=���1>��]ܡ�QMB�g�^l���0�}l���ޤa62�N}���i`��>��T��$f\۴�6�0h>�Y*��
]��2.�3��9��EK����}��H���V}ܽ;�f��r$�.�E1.qP�ENN"���}�eKSy����y�C�N#Z
�uٶ���ZC��I#����6���66�E))�Q�.��"�uC��YϨ(6.6Y��!���Β����ڳ?IR��&�q�A2������2�jO�K\в�0O)�3�djW�I��KmJ7�k�'�����g#���ٜ�������]U�Rd8��bM�P�=*2j�l�jMQ�kT4�:ٲ?H!m�KӖ���2]�:�J4;�����?���@_����jJ㦔���j�5R��;���&���*^
o�g
�Z�U�d51<��"��t�?� d�FX__���#IL��e���v�O�s�;m����ʺ��.,w��g��s����P�C<����u�-�k�%A�������N��+�������)/]�5cG�or�K��p���z�NϮ��f\�>��-����_;�i:��g�N��i� o47)��������d�_��7'x�-��9����'�Viy�S�&,����B�^7�_2�ӌ3ߧ��l㛕B���.�\�&#J؎�� ۉ�o�k�4s�?q;;���'/*��FeoX�I#��<��]#�|c��s����W�����������)��O���C��}~��C�[�dR�oZ���'����.b�#�T�_¯���d��"����������譩���l6sܿ�H��"J7�Io$Ͻ��6�9:z��]�?:ƽ{%n�XQ���X�[�2@[o�h��\%������i5�sS!xҍ��$���U���y2��i_�V[{k�/_��W�Ʋ).񞾉۷���&��;���|Af��B�1��uyme�p�5t|��v|<����%	v�����I�ԣb.N�&P]�;�Yu����P��I���'�{�K-�^��d,l��ݼyG�ז�\>#�������4J+k�2V���H��һP��߱�TE,Z�ӈkX�Qvߓ��{w�tS��TX�!,��.�>h��c?]hL�e��-{��N��i�{�1����@ߢ��6�e��5������������X�����D��7�ٹ�[&8�/�UӦl51)��ZCl���w��b��t.^�ԑ�\��B۞ks*�?.F38;�bB3�PT�pV��'mhV�B�jZZq)�DfC
Mna\
�'C���l��pU�B�%Y�����TZ�+Z�m�jNp2�-�]�G�M[�a��x���|����l���wxBE֐>�<�oU�g��	?/���4s3���l��w<�M�v2-K�n����)��
�� Λ}��h�
u� :Ky�M�ϔ7��@<4���+��]���~�%���T�j�:�!.u�:W�@�[�'����0&���[	V�Inܸ�����^#��H�����Mf%��:�Cĥ_���OC�s,�X���0��!3��ɶ^����_��#��>^�D��|�	���v�6w��AWh��ԟi[h�s\!c^�6���Ks\�s4�FC�i�X���&h,��J�n��X����d���J��3<&�;�844n|{,�~�u��v����O�̾�?�')3k�ǖ|��ʸ�	��eS��u�,�B�b��4�F�]P�ik~I"ES~rZ�����QY�4���%��[�§R\����w�����F>�\/�g�/�ެW�49���[�VU���}�g�p���H���C�/ta0|g���|�+^����(�")�Ù!�9����:����x"����t��� �3��:�[2�%�'"�x�?gt[�����˻߻C��h�����@�f�E�?_�&���A�m��N ��m��󺆶<�z�BoXH<|Ȃ�$�|Qђ�M�*6��CL�����]%]�]���kJxcV�zr�a�}%-���<�%�5ۧ�K�]1�4�r�ޱ=��U�b#<�(�O!������(*��R�����S�OC稴� eW�B��^;������` �'�'��1��ۡ�D3t��5�� ��ӫ2�Wg�q�Ү3]���3��T�U�LO���
��`�Q�%�֍h^���{�6wiq~��gT��
Z��G�e�V���dCw_>P�����\.6��OL����X��DE\�T���M#�G�Vd2�/PnEh����Pa=��p�7�;�x�Sƨ��"�L%)�>��v�X��� �v*ڿ�ͭ��M���!UYT��׸w�)��� ��Ȣ0m�(P����'�=��ӏ�>~�gF��+���ё��*�W����)�v~[�oȿ�y�9�үv�\kU� d/���Z���i�1��_����	����� �y��i�	���.H"yO��\�d�oZA��_h��#oX�@���;��<���F��jqx���_���|z�&�7��{���<S�^I��zE߇{�}ݻ7b�?f�0���)]�G-CF?�˷��c��׈~��iqr��]����*?��<�<����e��O(G? τ�$����l�]��|*�{I=H�C�*5{���⚛˖_��/��*��Z�Ũ�}�k�a!������9��xSi.A�u$q�:W��F�\z!��sĢH+ݪ��I�Ⱦ*��7c25��JO��	m �DR=6�MD~d1_I����x���	%�Uh�������6*�Uz��ʸ��;�O���<��������p��o���p
���N��`�"��F|��8�`�� 6N�����-2��2�Vw}��4e��H#�=3�!�5ڜ�Kg��L�B�ٌ����oR9{*Fjr�%ڛ�;��(�>��{{����
t��\�J��e�h>]����<�O��ݹq�.Ѐ��A)a�[�	�g@mC��-8��"�����'(No>��\IX�!��N�d��/�~E00H����iI�{�i��v��c���1��s���k�xf�c�>n�]�Ů����Ռ����e��dN���!i�hx!�֝Q$MB
^�g+E qx&�)�M> la�x�1�LT�vɟ]����j��
�!=;z����@۰�M��Bh���*q9��*03N�~I�l�gK4@�����F���:��r�c;�6k�~~���7�������Ü�4Y
Լ�Y�I��v��M�����+4��Hm�:}����o�KbL@���_<�AG�3j�(�=��z��N7�>�ɠ�oh�Wfl��z��ɏр���_~��_�Dп>O-�%8d>����._���){�l��G�{��|j�ˈ�L�&���+�pD�^���-�P�!o|��G�.���L� �/����`��{�Uz;��3wmq("DP�!�l:%M	%R�:�XY���_����I�<ΨGRB��06(�������m��d�|�e��>���[��/1{�`�xQ�<�?$-C�Y���Iǹb��lx/pR��j��4R�)��Q�������DM1���R zx�<V�N���1N|���O��w�����fu[���@b�H�����x�{
�=�
�����+��JM+������
��g�QC�>���׽K~��N��ɓy���L�����m���e�ҍN(O�(�yK��W��q��湂�`[�f`J":do�����2�Wg��B�|*z>�J�U)Ӳe���_����N�����o _�_%�ǧ�����hD|v!��;9%�ψ=_�i��z�艠��UYֆRE"��� �֗x�./�ӳ����g^�����>��ۈ�)��ڤ���TDgG��A��6AP��á�l�I �𕭃���oO{���cF��|�Q@�w���D6�T}�d��ޕ&ɀx������Ϝ��+��1�	�!>C��.�0���Ҋ�j+�����s��7��,}����R�8)�Q�+��<MM��?���>��;I���K�nӝٚ><�ݗ��TF�0���k�L/���裏$�7��U���'�Oh	=x��Flt.Ni�xE?���j~����?�o�=FI>��~T)�#RԆ�{�ާ���{�"%��W��8��֎�c���|��7�F��P�aX�������kjZ�U��j�#����;c�I�R����5Y���X��e�e��	*?�ZB�"dy%q��ݒ>�����|,��D���P��tqc�`g2���Z�ha�9 ����+��QO��$�����I�G5j!�G���З(����Q�T�*Mc�kѱ�����H#"_Z�VY_�ȧ�J�1�|2�܈���!��u�z����ڥ*z���6�v 6�P�!�B|ðY��a�� g8��w�1�������j�T�|A5����ʌ>�`�"EG�]¨x�<盏�!ps�N>���˿F{�t��1-7|r�˞���(��;u��iF�fE�{���}�����v^�AFF��G���I��Aî�tE��?` P�x-Ǵs��`ßՠi:c����3��w�7��8��ђ]����-F)'s� 1"���$�{F������A����� ,��Qa�4c:�5����kX����7l%�(a_���R܄��������X'oJ�UHFY�G�~2^у�L���ꉔyD�%xFQ{_b����i*잇{4	�7(Z�&���^K�b��)�c�K@_�ߣּ0�z��A�
̃*,�Ud1�s��H$b�>Ak�sF7<�#�<�`��k�Td+2L�g��D��;_�����-�?H���<����cF�������mس+�{"z����f<'��9�a���S��	[�����O��7)�M��w�	�z��Ox	~V�/�s��"z��*�7�nMP^=��k��D���D_yuD�?፝]���3z�lC�Spkv�w�]z̞«�|��x�~��,ۣ=�RT}����> *���f�v�C=��7�+-j���ݰ��$���~L�z�q~���(V�O���)�8�E�>���'�!C{?;qB,"4��ؽ�R���UǠ�����;��w��1�^?�3���y����;��%i�����W��p�ײ��=ɞO�̭l��f
�)�8B��%�:rcNJbH M��#�\���'���z�t}b�
���.qb2h���b�C�`�@hC+�P�y|���ZK� �תQ)�(�Uy�������F]�g�0؛h��,;g;Ȁv�N�kc�a�^�x��|9��[�_�i�w�Jկv�cOi	��F}����lv��T_��wZ��]�V��:�v͒OC ��aNΆ�e��E��{-+'**ٜf�� jwт�G?�	}���ӷَ#V���Vz���}޴o����k�G�A a�M��¡Z�l�Z�$j�#8ɣ�T<��5��SE��`lj{sy<�͛T��7�V�N&@<3�'R�L�&;1�3a��w���� �%=��ic���	D�ǃ�� I�� �U�x�B�uc}S�l�J壝�	D����R`��ā\h@�C��Q�*�#�K�������0)�ɠJ�H��r���$��}��R�t��Ε!��;��0;�
���������>������}r���!��>�u��nؐ"�2����o�}��!��o.�͟'����D�/��~�]:z�b�����#��y���熷��={��k��"��[�ՙ֝���_�}��:/������=������M��o��������D1�J�9/N��B��FrI0N����ȁ�X
o��:����M`o'�,�:$�M�W�g�ڌ��B,����qU�^���1��f.�䠁�I*�Z���V��d<.� ڡǏ.h��w�z �^׋� �z��;�y�i�]�Œ�U�*�_�"�-�J}�|��##t������T2!���! ( }Q�$]G)N��B�^/�5�Z�]p��z"y^|&޻ ��"*q~6�A��d�<zT�?�XdC�=T�R�+������G���57�q�b���|#�Ic��/��Z����:1"[?�uyHk>��Ha'|�)e����3��0�ϲ#zz���o��X:$}�AFK�I�Δ���w�1�`�um?�?�,������ҽ��hq�<>q'�a��OhroJ_������ɜDnSk'I�Rx���=e�<����?��uFS��&��=�(*�vyA�8�WK�j���,F��5��<a�Wƅ� �ڄ�?΅�qo�jo�c��*PU�u�n$��֔l2�y�j�!�����Ot��ri�������oz7eD��p���p0%�<@S*�@���G(hxW 4���kR����Л1�9{5k�"��9�=f��?�M j�g�&�U~�.��Q��(��A�>���������T4����w��N������qM<$��_��<H�b�c���嵱��
�o��M�Bӯ���<P�2\{p����]�~��+;T|B'����<�[�u*T�(}�r���z���YB�t�̈́-�)�}-���_ݠ?xo!�R������+�Χү�v@O٠���R�p`Y �p0Ѿ�;|���F�wP�"#F�?f�&�c4.���:#{��򕄶H0{#��;�R���u���}3�4X)�6l����y���2�z��;fT^�ƗDj�Q=P�)�ߣHy�t��H�`�q-51���5�̯����IiV�l�.i)���W@��ɹ�IA�y�څ�|��L,����Lm�t�(UW����ۀ�.�o<��|����
u(�@�z�i��O�� M�#��^��4O����vR���̄�vZ�h�`H���1惃=�f�I%r�;"3�q�2��
}��ȗH.�!P�A^��ܢ:H��T_���ɟ�zs�"�,@��/TbṪ�a�V��y�QԲd��]�Lc�rC@�VV��ii� '7�������)�����������*ޜE�K����/��\��_�	�Y�fZ�&������h���|�m������Lkz�[�_�����=�BU��Xb����j��|��������b���&�ut���[״�Ç?�r����"ǱK9�3Ε�"��X��_[�>Y��R�5�@<�(0�)��ѣϿw9aX��*�/ڪK�\�^��.��t���(E�Y��</��k/(�A�26 eś(o㪉Ur#�P>��tV���B��N�{���
3����=�nK����ߥ��,G�Z]��!)��_9���G��_�K���D�q����?�u�jN~��B.����׼Y��O�a4^Гcx�K:?_�W�1䵱�_��C�:��ވ��鐍R6�$q�m�шf��ӆ��Z�8�bg��אFa�=)5=���xb����k��v;W�����<7�L`͏��P}W��ilEדﴀ4��5�U;kn&��6���b��k��[o����x/b\\�`��d|GĆ!G�Y3z\>푀�����4�P6���$i��
M땠��p0�7��Ts��)��Vӆ�2���,�_�5:��"4�+�|�{�\	�Z�LL��)�=���y���l/�����?_rk#�?�����Ǡ�f�.�u,�r�x�h朖��V�́4RX�?����'C�§�����Ё�=L��Dc*�%],�������	�y����	%����sC�輤ǏWtm=oG� Ľd�����g���x����96��ʇy���g��
��*oT�l���{�2t1;�D��ޤ�3^����7}z~}�#�=�&w��Դ�ײ����3�y��:mv?�O'��w!j1ǚQC�!At �O��_I뽈��3H�=?ƭ������R��M�5�]��==8��^w����j(I��T���������XҐ�s��`-�'_5\x�T���hH~��	�2+dq.�RV�������0���
�9
�He��|���ċyC;EL��&c6T#��|�����d��g��?�CQ\A3~-d�@}�z��<.���ޝz/��d+���y���C:�M��կ]N�?�M�?zN�#��9�]�:�g~/$v��m�A*%!\�>M����{cu�	�GD�B_����O���)<ƿXIbT_����K�E^�_}�u��A��}<���F�:z��f�͵����-_H���($���Y��Y�I����F<�r�Zc�	n��	yְ�i�O?�t��Õ�j�,�6#)�V�3y�s/)�%�@��J+��=�����0�ַ_�*-x����M��"	Jc���P%)�=����Q �$�%�jQWˬnZC.�,����ݠF��9xW�{ ��ɻ�K�?��7P��F�m��-�Ӊ5t�FS#�e-�� �	�:q	%���[o�O;8�v����*�21X+��ß_��W�P�7��w��My/��5��JQ.�J��'Ԛ����l!��%r_������ߤ��=�8.ħ�B�dR��o���E��Ĵ<eP��Ӂ_륰����i%���^�x�'H�4�Jcbp��>B'�����_{���B�𧄐�4,g��"+�?4��Xk

�B��#n�{�D߹s$���f���>�sd#��S0AVb��9�YL(������+��#�D�@�;��HB�f���pi�%QK5 �tW�P��}!��\�T��E�!S)D[�u(O�`�1��'����	���"_���(1^�\i�ɷU���wqb�j��O$��R�\�K�s_��.������s뭠���^JhOdB���/bx��~����xM�p��*R��U�=�h]2�൷ˇ=ܓ�����o��N� �g9"Z�!�M����"3�M�d�gԠB�V��k �_��j�W�T�����7}z�=�{�nIp��?]g�'����5}��{�t�����r����~�4���۲pm��o��v��Xڴ��p9OM������uo�ƿW�DM�H�(ո�/���'�{D"����E*�A���H��Çe��^��J~��kS˴å8���q��7@'���F`�UmTY/Uk��]���zQ9�"i(�ּ�����n��kؖl�U;��H��{��_!w��X�kn�tJ�Z�UZ׮?$������aP"��~P(��¸�	�C�j�R
�*�+��7�mvq��ή:�A!o:��b�|�O{lDnܾC��S~�'�Uש�4حE�0#��{
5 ,�Z�N��yFg�p��F�w��n���;�O��q�T��6s�a���KJ/�~��F�w(J$�-
z>�p^<[�{8��?őO��}v9iAwy���1B(O&��W�fsB���ɗ�}9A���=�C^����&#�{�+��z�c�C�����E%,�!*I�5
Jx�&���u���_9do�6��Y�6�ٹ��c/&B<}O��
B�fV����d��.�_Kا6�������S.bX)�D��lT{J_e�"�o�68�H�Nw�P#F�^@Ii{&9�A���l�Кd=)i6�a!��`�И��� �V4�<�����;;�AbP��O�d���W�����T'�{v}*�x�o��lA��#jf+A�4�o��^y��_�~q[r�����JW��t����-x=}��k)���~c'��[J�8a�%����|B�g��c�>?���\l�O�zE�Q����ʫ����=։'r��P�$dK?��!:�߰����V+��qJӾ��m<�P�,�z<���y���#�:c��)Ⱥ�4��\�<a0�q/M�|s�Ƒx��r���Ƅ�4D���V��f����?�1=��nA8P���(�V�
(:[��;���q�:�?��ZT��x�4.��&�~���k<E������{�o�`p�A�y���!��4�Ǐ� J!�<��op�`�v4�`'�A�9�ӻ��3��|��EIg<��0�h��?�=9��0;t��^#���=G��	��.���Q��8������3��R���Ь;��C����d.Hի�H�r�QX�<��R�i���hRB��� ��g4N�iww@����l�j��]0T4_�6�dOc��]'��h!���0��l������ l�G�o�A��̵��T��uF��x����E$͒��o���J8�@��E߿Gx����Ь%W��Ĵ8Is�:�d|bz!���E��i���ڑ����]�;�Q��3��S�.�2Pх0 ��6Q���{�V:")�ĹVR����@�����oH���m
��R�1�nɡ�=�Q(�+�����X���W͓2��@�\�!B*����M�>���C[5�`���GҲ��,�#7�:���!�z�<������	-�(L�(�Yr摧U��Hc���j9����ƽCH}h�cܠ�Ci��֋n}#��V*�'hʰ�A+O)tu���I�EV���U\]�������� ���ᅵ��fU-^k(����Wο�礊��U5-Ү���[睊=���p�8�:��IS�k�q�<��D_Y�z?;=xP}	�(�'pV���[��?9���T� 6�u�[�%�<	��ԓѰ/���̰��_��qI��W!�����~�����D�>	� �k��c(������zU�A� �Dȩ��n5)��Hn�7[�j�0�|p,ό�k���ZM�?�x({��"f�`�9��]��
�+3�g��6-1����ϋw�?�'����}�}Fk7���KF�7x���
��'h3�Ilk���_��g��f4e�t�6Q�J才{_a�r]g"�|v��m��)P�jƈ�7�� hi=ȳ�/���4b�S����#���R�~��OF��{kz�����x��ɞE�(̋m��n9tý��oB�7�t���^�K8���1�K|�����]f���������@\�R*+y�^<�M�(i�F:C��3���I����|?:r1j�_��R�j_����� 
�<�&aA�S����
C�x�������!��f���&���^{n�-S���Ĉ��J4p\����x#�°��C�&V����G�*ל��=g��K| .:�Eg˂f����#4O�t��љjʮ�x���5�<��Wͽag��$�,y�A�4�B�����u��0�P���(J�{d��<ͩ(FB& ��e����&8I�!��6�o�w&���Ih��h���W�HF�0~�a,bkr�׹ƶ�C��Ȍ�i��BE���5;�� k�M��ǌ��Ψ�D&F�Ck>��I��BR{ݓxn.����u�jB`�r��]^I�AP�dj�"3;=M[�.�Sy�Ua�x�QS#��6vC~`밑��3 (	�H�uF�nÍ�Z����0��kA%�jt1�$�EZ$� b�����F�yC�G ���ӂAN=:�^Hm�7�u1��J�=۴盗���Y��v�紖NlJ���-1X:)��]v�axN�������%]�"[}eF�7������r�;��K�Ϭ��7b�)�8/2sM�L��Ő)h�}�(��W͚O��kU#���~����E]�k�d��̵f��|ؐQ�{8<,(Y���i��o�C��hv#�)H�*I�ڡ��J�'O����D-�3vK+3�{`�G�J8�s��*ʚ��%af�L?��Q���Z�����77�,�͈�ea��-�M6�<���$.�E����t��$i�{Q/nI$����Ih{oP��ue��V�=�HF?
���|�sX߂��AJ{;4B��k�7*�A�dt�|�*\mc�!���$z��O*�y�geLS=l�7yk�$��ɵ�ulQ�a1L�s�NC��d�1��Hi'S+��K�����O@�J�䣏fBa�J�R�7eHh��u���.�ޘ��:��n�|���G�.�L� 0`���Z(��a�&�
��N�7��,+M�,j�t�"�.9(b��<�ɯVcErO���+8t/U}�u�ZA�.�\^zn{��:��V��Yݡ�{��CG����%��2y�ᭃv=�%V��q-c�3�g�K���� �Z�~z~*�-[�)e[�^�	�)���:��=Ĥو������\���ʮ+3�����������,6I��.7��\2� �1��"�̣4Lv��ky��C#�3a}���o��rV�C�;7�4�Ź��|4��/�@�n��(`#J�<�M#��%s?Z�['r	����1=�A�~Aw��4��pu紷�Srm��o�.|����'��r�,\%��M&l@����$W��P��(顃z
K�K�a���P*��"/�X��,ll�*��Z�WH�#g��{m���`�j�HSmE:N��:a'���j[�Z� �1�t�����(��po[�y�w��R��"��}��G�f�1ڼ���_ƛr�j� L����0U�94�V�*�V(�	��6j*t%*Գq��r=J!���H�n-sOz,h�Y$s���ؐIG���s?�^�X��$E{�]�N>�I?�|�������L�,�o~�^����	��*�Q���P:��SA�5�ְA>^v�|��2��Vabm�ݜyu�����0��U��C�m�l��q�&�(�6O(��x��[�a[ <�:��!_х9t��L�HVf��ڈ �6 �4�[6��ݻ�'��)�#��vSG�%kUas��/��m����ɧ���x+{��AC�bxA�>�p۟�
m���1�t
�����9H���y�hp����SJ�cڋ�SGB/��\���1����v�����w���q\x W_�E�^�p�ҕ�^=���^��R��� O�]3;Y���+*Z);_)%ngL�R����^b�=����/��ؠ(HB�3M8J��◎_�Io<����$q�_�L�.�-.�e���&�P!\���(o�j��!@�ܼA+²����cO�M�nir@6�N�}��,j��5�m��}�(�� D�k3��z�zl��כ#�Iܿ��%dS�g;���C�!q��>��6/Bz&�L ޑTgtv���3�.�1L��fn5�((W�7S�<��DA�<�:�Ё�&4��"��5*h�T��a�����%��w^mF%rF1c'2���1-kԄ���[�� x�g��0E(�s��`m�]��BK�{Ì�oU����̶tu���?�`����Ɵ��v)9�$��H���1���xd�Gr@��k�6�U��Q[�?wp=���'9��W���7��[����q��d�O_�*�������z��'@v���~x��?��Ĭa^�%��m�}Q�	b�@�e�����h#��O@#��$�T��7J��'�9}��g��?�7_M䱭��\o �&h.�����R�_�>UՎ�#qY5 �w�hM�ʐ�A�o��Yy��#F���+���ʌ9m5�>}&��T�G��w��浩T~.gs�L٥�&���y��! �rH�<Tw�+�47�3�IOF�l`(Tb��ݰ�|V���l�&`���W?b�(hZ�e*��#�Q�
)�Yi(F	��)�_�MN��ܦEsL�R$$�/敢ݕ�Xq�^3:�+�1�`]j�1f���J�G�^|WHU��6�
s�"n�K=N�A?��6�@s?��.��`A�Բ�5����A�(��*$�BJ�$j�F�Y�ZH�(=8X7`S�8>��m���%y� GI,�*�Ql��-<Ply*��	����kThz*�jB=���n�˃.�Ś%�"����= -7fl�1��Ib3a�7���!�-�	m��'QƷwt��u����W�[�p�y��8b2���=��f;L�Υ�g�uFWM��if�j��s`�C�5�Vx%sl�']�6��ɟZd��&��IM���0S��_��1t<� �R����~qxns3�w��C=�2����F�EAPm��n��(��jl��	q���7�L;�?~���V*��*�vЉ傜b~�m_WB���Bg/> ����
�nd/�.^�#��S>���O�kl���R������U\Wj��;�P$.���D^.�ж�q�$6Wn�J�Ps���5����h�;��=�^s:?׮>@;;�4�@3�Go|�w�#�8��kH�$7zҞ�b���@�f��A���Fr	��,N���8RjWΈ	��@���SiR�X�4�B����hƨe֝�+F*�)A3����Bb������}e6�^k�4�X�q[����1N&��m��-ߺ�*��� �p;׾�f;%E�WM�9=�n���
�@�H�	�Y�� �.dd��06�C���.T�o=�3�z����별��߽�g��7v6��;��Gj����G���_C����t�D�#�����5ݺU��xn�B�CE��\��=�V��s���}7����׍�cE�g�Bv���u^��g㖛g�E��I��v�u]�5�H���S�Ϸo����x�=E}}Ἵ�"�#���_K� ^�k<���=x�U��!�0Wf��kJ{�z�箞�S�4�*�hdO}��C�^c���<�d����=D��k�{3,����9�Sd�,E�~�ԁ,�E`ا�XceԪ*
� X~�'�Ѓ�݁�*��T_����SL�٨^+yB�<a%�]�t1�H�z��<�L*0I� H~�ٽ,�T}�_N��ܛ����*n8�."HP���bNG34N���k ��Kr����&�s�3f�9�E�'d�.,���*��EE����KȖ��I�,�|*Ǟ�[r$�RQ�S�]I~b�F_4i��O&F�Z��=���h�� @�!����lʶ���:��sQ�L��4wV�I�H���l�X$P�Fa�Ò�[��$W?f/ﭝ��p�'ǀ�[��V@]��v\WB�3�B�vX��iQ����G�aH�6�4���2!<��
ʠ!����o�JT�F6{��ZF��;	���P��q�Y�&�$F��U��ϲP��ڌgc�P��
��q����B_M�c���+aĔ�v;�&��pE�ꈒ��������-�Oh4�5��z	�^ߌr/4�l3��G����ӽ�7����qYn*:��xv]�Q-E��1�I]'�.k��ʚq�����31�yL]�^�+��Z��v��,�̸;I�������<v�{�1��k.�[��QBMR�.򥴁��yd�QP��~��d�{��-�.�a�h2,h��i'494 *ϡ���T�X�%ۙ����#U��~����F���
�P��6���i��_�ޣ?���K�87��L�˕�cKh[�8&���8��z�<8���sY�������x*�^�r(4���NЈ=-h8��3���~+�F)�q{ոb啘��3�E����'t��3�3���\����<H��wJZ/��	�4Mw��E1�H��W��&�$ ��PEr �ު5Ʋy� ���36�q��kF�pǁ��5=�.�����r/��tn���r��>W�)���0j��� �8�*}[���m���'5A*�0���Z+�� �̬�N"�)	DՃBk��R(���=�����Pf��eqI���k��h���gV�A,M���P�{!/-= ���%�'�� C���B�=�����ۜ��2 Bq
��@���ޗy�6����{�����HLGT6���E��Ub#G����<T��׎�Xk~�r���7R�8t$4gt�iՅ��c�Y��Z[��)t�r^a㹼Td����5�Đ��o���֯K̺gA�t�VsA���P;�\�/.�4#�IY���K����0VT;��4���K�4�H�)i�?_�
8�\ٛJ��jH}z�ؾU���\a<_Ƅ��Z�1Z�4�bSк�������>��y�#7脅$�Jl߫&Ԭ7��_/�Y�ᰤ]�a�Ҫ%4؃3یD/#�tA�
:���������!e|mD��c�2ִc�ҽ��J;`�gs�q�����½�`I���E�4��E }w�#�*A=�v�����B/�� ���v�
���ٳ��\��i�Fd��F�X���U��v�^�K1[��#J�G٢��O�t\�z�t�A�ּ���� �56ɋm�K���CsB��M�R� �;6�����p���]݃ڰ�S5�".�+�v��j��^�\Щ_K"=����B/6sA�a�P"�ړJ�tYhZ�M�^/MY2���7���p�1J�Ċ�ЉЬ��ŔNOg43�ܛw���8~A7o�{t�����ZZm����7E����칬A�>_��Oi0ݥ���"!`��*0�)P�T�^� �w�m	5���C:/e� 7#��@=�i�C�Bf^Gi~"��5��[8/N����)��C����`q���5BC�n��k�u�W�6�	�^����LBsĚ��By4�؁��t�Yְ�p�%nc'I.��DJ��;���.��KW	��QVXLaK�u����\�0�q��x�4ǲ��/y���d���	������<_�W���	M����J%�%���z��'�<���'�X�fV��U]Wn��r��)�"ֹ��@��з�x�l%y���Z�饗^��_��]γ���-����
c�4��]�G2����z��B�.�!ڱ��M���)�UT�;���4 �M�^@"�ev��o���pc�`��D�
���d��T���ĳ`��3k�햕G܍�+�Q�OТ�V�V�rYu�\^뾻�eFN���ם�J���&#�:ʦc�8���ƃϱ�ￜ�u�sy�LBF>9-\?�60\�'���H�.X/�:K��Yl�����i��b oݺ%;F�F�	�GQ(K���v<�<H. Z��y%����uS��}��Mz	�-0�q$ެ��D-|ބ���(�9��9
��f��%c���Қ=�_�F`})N��Z�QaD/���*Y�Ϸ8sd��1�ԣ��R�m��|��;v9)�J,no�{ʴ�m�y���w)�O��y�{���m���Ԇq�ɵ�l]J�^�#�]?�ݛ����Ol�A {%J�	�����b;J<��y���*%�R"�l	}���sL@*pو��g�R��)b܁0{��W&ݺ�&���J���@j7~�~�:=x�]�0X;����_���ݕ��+7��3/D�U$<�OC����n�2��?�z���c�q.$�P�"�uʧ�c6��P1��ݾ��/,BZ̖�ٳ:z�::�Z�b��>�u�#f;ldl|�M��Z1j?yq!��e-��B�:�k�����}�M"]ăC>����*��$e5�STC�
�0G*�[*-5`C�;����LL�O�L�c�z���l�s��e�59���q�KRʉ�y��
����:���mV��h��v(K��Kߴ��.6�g���f�����d]qW�c��A���B��-6&�I�<�#><�{��K�Fm:9�(ءw�j1�~pAI���8@��!���m�YJ�~w<6�/�>(�Ewh�W0�~^ĭA�*��MJK�\�w��w�oo�:e�����#g;<I%2�9��e�I<:�4*3Kv�jT�5��:�5�2
��¹X�:+G��JBO�*��H[�F���Q*a�8>��S���lr�0�6+�DF��C�Fh!��)!Xn�]B�QAi�z�h7��h-@Z�YO�6�X+���W-�����sg�Z<:�D.�un�[�ʊ�pxe�~�~�����P��z����7Jx��������-�"8XK�B�]�|�I�k�V��@n�C�2=��9��7����\�&��oiC
Hz�|`¥Tt�~M���]z��f5��w���/��Wr]����/�S����g�b��۽3����,�ďC�b�U�D�B{0B�lH�t�ZP~qA��TP�t
Dğ��ͨSɞD��?Ռ��}�ݧ!�9 ��߬|�?�i1/h~����Pu�o��Qd6�{W�9��d�$���.	�oem4�r�=ߴm�V1BF���e�M��BY�zk�M�M;vbx<�T&@;�4�e͡��bQᐸ!�6�y��/'t��^��Ȥ}�Nf����R��o�q�q��<��N�6��W�%���I~h�j��K���I�@����D/�AQɆTs:��/�EN7˗|�&tx�MG)=��Z�U�Έ7^k�5�B�",Z�)3F�b�lղ�ܳ!���̒���h��x�$i�����ǭFM���z�Z؅ͷ&~^���FK�U=��< ���:�Z�A4��r�!���5���j��d)\xK�����_��4Y��`����Ǣ�\r8�ĳ��&'F%v�w$��p�`kT�*x�G���N�Ǌ�RW�ꭄ�o�������5Nmn,P-;��4Ȣ�$�m�3�
м�39:��~��r=���z�ʗ�؋�+p���Z~�����E|䛖=��]Wn�qy9dZay
����7���M������BF�@,)tx�5�M���g���hs2�.�詹<��h0�?�d<���待�rv�	��hu�^����R]#��5MP@�y��p��Bb|>��cFf���:YJ�Fy��skT�)��Q*EP���(ʗ�������c#qϊ�o�p��\B?<�PKh×�>��\�K���n 1�2�>�K��2X��Z	��wZ�N����^�
S���84b�E��aj�y Rd&%!�ch٫�jH�-�kף+pQ�+������9�={}����f?Ƚ<��zɇ�/�OP�uo�X|�Y�j%ݓ�J���$U�	��d��U�Lx0�C$h+�`ܠi��a����B!ސ�kHD�0�*Dy�:�NJA�+F��v=�xJ�ώf|�L��}�����$���7��u���0�B�W$��@לl��B=��9#;�F�؅d|�@��$#_���w	Q�VZf��!đ�L����x���Ue�=z�C/2�|���#��.z�6�ȁ�jy�v��T!��L���2�X���;4@�,��I�D諾Q)CBFÅF4�Ӱ�������������ڮ�=6 &O@�Av�
�=L4'�5"R04D�x2U�����Ju#�=���c|�PE������|8����^~��~R>��N�
��tҗp�c����4����*Q��1?;�����\,x媚iF�7���A/c6��[ �%�D{��t�	�'�͋�EG��q�NNh�>��2�?�
79ζ�4ފÛU�D�]ɗ�@����Vջ�f��@�YY���D.�`<��n�oJ�KK����{�������{����tmBV��$�e8A����:�G}t�m`�s\��L����_﷑琂�00���(2�������|G��^��ހ� �\�"kxO�#�t:Qjj��ǷX��H�,�1z2�A(]�"�um�F|W�k�2C��t�p� F�*7����i�$\b����RE=��g�v��c�hUO�<?���Gep.5HU>���⌾{�Kb��C�U��r^������3OZ�}��8Nm��b�.Z��.�/�6Sau��B%X!�*����6���z�WrkW+��]V(u�\� ���$��~쪨����8��F�'���5�J��&��Bg�W�d�$n��@�B8.h�e�-�阎L��ٜ�Κ�E@����\_��GUi�f�Y#�e��<�������c�}>�So0
��d�ٓĂ��'��{ʃ4�4��f1�~r*j|?��39��P@d�������2��g5%l<�s� l��6&����I���`��f���]���@� }���eA��b��fW��U(�rON�:��n(G	��x@)�6?>���v�B�_��z E��"OE�S� ��B�n;���%�H��D�F蕈 ��\Z�q�q��Z�ՙ�h}�lTu��K=�t�mu��:��AE��7����C@.��׋���3��8��
�\T4��c1>�r�J��ʐӔ����=I��A"���v?�~��xgf��.VmvAuf�eC���-�G��6_��3QE�*ۀ0�H7��d�o��$i����������Z���B�"$!��H5��7�'��<H�z����u�䋗Q�����^2t�zW�P��Q�:Pyjx� ��V���"\���5v ��� 2�]js�ؒ�USu�U�Dʵ;4#q�h�8��4-pAΤʫ���D�Ȑ��	���-'���oVv�;��0�Y�k!Z��c��+][Q"��B���!�������Fx�I�@���^Y�虍z h����Њa�����1����6�A���C��Oh���c�ǋ}�nĴʻ�U\_��W����d<h��;��K�W���c��<nH����ق�"�A֎S��h7��g/���Nz�*�=�$)F�MZ([���|A;�P���/�(�
I�N��W.Ds'M�Td�l�ĵ7��Ơ�!%��+\��,l����	�B³,�J>��xx�����0�'���[���&�7$�F�|q�Cc�=������3j܅�l
�5^%��6o5�>��y�Q����\����{]lZ�x�V�E��/@��ź���$���|�F� �x���E�	E� �,��#>8S�c
�-�?�����:1�lU;ݝ��*p fhi��$�ʯf	�T��U� �2)b�}!|�<^y��ǀo�*����M܎-�� M,�c1�Du���|#I�M�s�x���Tg���o�]s6��� ����]\�u�rAa�܋���x}aF^�K��wy���K6:_���y>�ϋ��Ia$��3T�n�釰[�I+�!��7�j �R���V"+D��y��U�ǚ,k��Y��x��Q�*��P����s�H���6���O�!�am8fC��+��֩�������x�@�U]_��/��j�b�=�¿F���ϡķv��Bѝ��邑2�Z�合ElHe���oS9	i]�y#Fݛ�L�jI3�۷� �-ʯ�ӟ��D�&��<Fp��Ͻ���,�+1�)7/�œ���:Hɚ��Y�݊a�5������h���K�B�>�ؓlȷ�+W����QԚ8��U��%���"��2(����Kr��M[!r�������;�u�z�|r�|dH���=�j�����!r�l�/�~�࢓!��Y���F~i�-��b����#��������r�z�H����U����4F4[n���{|�����Ph7>�4������PQ	J��@�LQ�5��
B,Eh�*30�ꊃ�GʺH��������J0�P�l�7��eUDDzs�ӏ�y|f&�������f,�"�xZe�lu,y�&��Vﰋ����z�28:J�� ��q*9	 mT�Et|�N'm�\B�@诱ܵ��\+̢0�4r0��P�RC6��Xh�g� G���X.�A�Sռ^�<r �,�������V�³�P�f��fp8���]��AA⠬Մy�TH����$6^]������HRc2A��Դ�q�Gci��K�8.���0���Z�	A��Z/R{��!@t"\�:9⨠'v	v����m���'R4y|��{<|�;|.�L�S%$�b��za���ڬ/��:6�䀄����h#�]T����[���$�	=
Z2�h���֟褅�T��rMx��Fn�4Aꉈd�$�<5�p�1��!4�CJ�ro#���BG��?��{�e�a��B~U����Y��Ӭ��29d"�r�	n����סRf.[=��8��t�{�;6n��A�G=���DZ �������:�x0+p��+�g�V�F�[إeՆ�l������	97�QI=���;ʦGFC-;	N+�3��+���XlC5"��m�2i�Lg�?v���ytS*E~��s�Ԣ����"ݲ����&Х\�3�X�2���R�Ш��H2XT����yd�S賛�����c�xmn�ӮN^�B�W[�n9W��wkX���^7}/��a��՗YptW���h��ԗƴ���
fC��2�_s?-#���|������d^�����)��*� 6Q��pX��U<���U�L�!3_]Ӹçi�څ���k{�m���H�ka̞�\kb4��)�^������I�ݨ8a�0�]s  E�i��k�24��[Ռ��$�Us~=���M~O!a�Pb�$�<T��#�|96Q*��x�����^�u��^��u��j�/�_�{nii��8���ɴj�X
b60�f�����"��i��N���K(!h�6yN������:40y�s>�/v4�R.�ݜ��/�%9�؍�n��Lj<��A�ං�FU�B��&C6�͒�^�a�@�6����-��'9j�37Z�*=K=CZT�V�o�Ո�H-H�����-��W����H1����f�k�?��y�H]r��W#R֥y!���ajT�X�oɒ����^���Ћ�Yx��T&��˅x�g��h����(aV��R�*r�si�����ţ��z��E7/x2��7 �4v�!:9���5t��2
r*D:#S5Jٕ��>`	�������g<��鿶n�W/<tO=��q�j��rڽ�u8(*Pv�%�ɳ�U����\$�#�(	/Ż1�g<,���l+����LZE�'� �/s^��L��U)�=O:����ޫ����љҷK]�Ǿ��.t��u����� Ђ���'��cG�9G�����h/�'�W:\H^R�Q1������������J�e���A����*����ۄ���.��5��#��Fk�7�fP�?�>��Q��$�CX�G;�ڠ��X�5�p���\*�.�����-VK�sg�ַ�@Uu��$ޮ �"���"Խ?�x<� ��JY/Μ_M�*]�9d^�Jc :Y�R�����F�6�u1���
R��xS�Gn��wF_6�qmO]��_U�,�{�4eڄ-?��e�4<OBS[F��;s���a�<�ޖ��ׯ9��pU����}���6/�B��`j�������3�k�k�Y+;�AkD�ǭ�6��tJ���R�׷K~��N\Ŭ�9��V଩�|
�ޘ�k-���_5߿ܽ�Ƶ��]���/�-�#;t.��t^\筸1����IƯڞ�K��2���L��$'O�k���X�k.}�ǽ�y/{:m>˒�8���(�g���b�"p�5�*$�,�~ !�M�w �+�|F�q#mI��a5DI)���!�D�#��RrH�@�c9!��q�!��Sa�T�v�D�ˎ�s��fDB��6F���+y��C>���҉�I �3؀�'���`u� '=`�[`?4� Ucb<^���h��`FM��Rml���υ���@�o��'�{��44�Y↖ᵭ�$��K�Y��n�{h�����U��.�+A�����Q�TWңO���@��?���P��kL�&�g��N��3�s|T9��HI�"��H�M�*e����R0�'�Z�#�O"*Kd���9�?Qe���*7޾�8��+�X��5y�l�N�B�cTw�ŝ|�� ��VX�G&�Beq(#&fD�|Me`A��,/�T����_.����g�ċ�IƋ��1�� ENM�rB= y>���'�|�u�z��N�AI������N��n���@��J���{M[q?DX5���$�9ʺ�GU��q���gVZ��1���B��"�Ŋ�yA�������m;t
����v#�g�@�<\ud�#p�Z�E86j���f�hAY�Od_z�?id.6�pN#�3�����Oiu��E��@<�����ߗ�]
��4�/���C1����O��D�ɩ*���t+��4m5eC�`�롋�i,'���c�\ʖ4]\�-X��`k4^���ژc�}_̚q��<"��_�⟮7A� ���������������iՂȥo��Rtf��:��,"�5�`L�k���ʵ"u��PcI�"�R5ʳC�Eۑ�̞E�i��<�M��6����J��yJ��x���5hk.��ξ�9T&Tf��a��i9�v<����hRjc����!%i�	8I���󺾜ѧV�]w��y���p���D֏���F��)�y��v]��}V-(�V�7�;��3��#�#�ˈ�]�!�y��mR���2��vw��r�r�ݦ���v<���*����;#����(�0�R^ߩHO�qpϢ��~h��s���6b��P<�Ƭ�G�p���f8P����1���F�O��h#����\ն7�{}9�M�|�&����:T�S���O<��5�*݇DZ#���z}xe,ȩ�usU�V�+NM�J�+递ѹ�6JF�A��I@��r%�;D�89 ����^�ě��чu�s[��Lu�p��(�6������Td�+����$��)pi5�~x֤X|ns��'.L���l�=�x�'6k���~L9�=15�u��̱�5&�U�M<5٩Ǆ��O���䐩>�/E����Ly��9�^~$��9�Q2���qDe~,��"��+�4���WF�� ١�X�L�Ф&xˍ��s����K��,��i��)�v(�]Π�ۼ�~���n�\��W��z�6�G�z����qb.D�7����tP���6�6w�.��^���K[Zl?\����d����^�.�>R׹�[�B�Pp]?�tܸ0r����������E�B��s��?��DU/{����2��~J1��} ��DdWd��~���H�~�c�璉�+=
������&})�3%��w�������!{��#���t��������R�����7���?5���G��t3 ����j�ΐy=w�s��ԗ��y��M긭���E�˱R����ߊ�:���崽x�>����X�lm��F@~�����i�T�����{y��}O���x�}$�߸n�u�D���|�9��V�$ݞ�؞-�%
�؃�F��H�
M�|�!7�_���Y��׀��Z��'�a˲�$���7��Ω�=�9o�]�A 3��C����n�����]c�b˳�l����t��w��x�燁�~��Sd������~<��}d�B �0�[�5���{F�YeS�Fe�n���'��s ��|����</��~���<�eR9�jߋ�����MǄr�Q�<}�X��޽�6&����q��	#��R��-�P	�7
��s�G�2�N]R�k���Dʇ��;h�H�aD� {�S�7���d�4%�Q������ *��K��X#C�9�!O�0�HM"�J���� ��=>�j��f;E?�E�	R��!^�D�e���q��S8Z�ע���wx4��W��'!��Q/�Ȇ���t��I�	\��$��qz,@��{��s_[E��kOO\¾�j#8[�y��	�6yE��_�z����F���-���M�w(�1���P#En�� w���m���"�!�;�T�֏��"��0*�P��1���Ï���#X|�w���%�����V���(�R�֍$m�5��{^X�ƺxP��c��!K��S_���q�i�)���$����-x���L��"���������@�־cE��'�5��蜹p����k\��R��r85u!���3��x��!�K��
��`�S �?���R'n��Z��5T��ۆ�(���+P�`kO������k*kgi����݋2	�o||^a�/q��HT��\v���8�[���D�Z�������5���g�]����\�NGC�ר}	%��9��a$��o P���3Z���Q!���q 
��\G��}㞩H�I�8����Cƀ$��x���՚�/������>�����w�h�象E���p�	b���!exl���ue��s?�t�����/�l�߮l�����>�Z������ђ��ߛ;����PY��_~���:�s���v�/#���녟ԍ��ם��;C�n���w??�J�F�[����3��X���,�o���.��v��k�������~X�o�l\��A�{�޽������ܼn���}^�˟��&���E��^�����X\���k�C߫�l��Cb�Gx�R��E��)׿D5~
P�	KQ�ש�n{:��jE2��z!��E�߁D..�Q��ؽǧuX(mON�R����+?��d�4���_Ht,��kF s~Պ�K�6t�+�Mǁ7{=4D��_�*Ա�����Z��3BF�^�BbЯ��7>|h1���D�.R]@�LJ��j��~�Zo�<��6=�2������ڽg{���y����?����&_f�x�qH͕���Z���Ib�q\��"\�@����c9J�Dr���-$HD���Ο>C6�D��=M�I�w�ޤ��S��D�j���%G���/��B�����3����W����3���$�z�mR�E4V��J�=�.O��;>�ܫ��F§�.`8m��sEy�mu�M~̎F�𡱃?�x<3�����ir�����beK���\kU������l��-��FBc� �^� !$�>`!0Ox$� �x�_<�^�BB�,�� 3������vw�>g�Z+��k}�Ȭ��{[���ջj9DFF|��l�N�_!�ދ�R���^�-�k����-�.W�`b����H�\��,����H�f���@3_�hM;pA1���uK^9V�rd@��M�!#q{V�j��؏1�	�V9�?�����1=�m�g��`a*��Bw���8ҥ����,�>�)�׾Ssl�Чr�wM�e��8���o�эj}��Н�2�����汦���ӷ����h.�7[��b�`�{��s���O6�!��ռ`nty@N~�]���^��é3����5���<\ÿ^%t���~�m�x?)�y��4Ȇ��]���{[d��/���m}-iDv�	��{Ά$� �3^J|�g � 9L�%���Y"PT��ڹ���\~ޫϞ��T�m	���)	Zo���5*��f^K���� �{�}�S\zG�yG�-���`�HH����d�˩��f��m��-i	cE��dSk����t��7�?'�OO�(�C���ɚ^:DU�%��(5]L�]�Cں�f�������d��Ь�ӥ a�8�Ǖ���5��	�$`S�!�a��oI��%�ͽ��D)?�<l�ߧ�SCs�����z�Q�{;yztv�IH�)2n�p
�%�7���X���yq:\e����q��q�8=@;jH�m�K1��=�M�v�E�'F�YO3�l�ߤ4�����gI0�/�z���M<O3�.�O�xWfs�<Ŏ�]�q,;��蔥M�b*��@q�6��2]�n)\V���^M)��Ok>��wD�����yI����y�i_�o��X߭�����M��h+�9R�����U�g�_�8H㡴^�B������4�l�'���Q�M3�<b�6���0,��@��YN�Lfȹ�qڠ��i��/�`��b7J]/�/��|�$7���h;�1L�8�e�Hֹ.����y>��"���^h/fz�Ag�m|Tׇ�r̥�N��%�(�Ik��894;��F��t�tө�J����F�����<6b����B8��M�[E�sd�U�Xjy{vҀC
E0y]��}}(��f���-�8[]�oc�)�^%D�ϔ��t@e�Yo����X�JE�l����l� ����2N����^X
Ѓ:8�NkFCj'�����7��dA���3��if~��l���M�WV�����!w���.�c�.������\/��=�m�<���������_��]��xm���l׷��U�u�����$��XJ�Zn�b]�����f:m;[<�f��}T�K/%ݚ�OQ��RR����z�N��	eEbCB���9"�n�3*�;9�NH�+�9[�W�=���0fqG�+$�}Q�0�ĺ���vݚ�|V$�!ۄ��iѩ݃0o�ͼ#��`��0h�d'�.���\�i�H�Lf�5:���.��n�j⼰��=X<�U�)��M���<Y�thH��l���}��h��-O��������� qR���x�.�6!��'�B�.�D�}L1O��3	@H\�Y�?�l�#J|��Paѧ5����ڙ"Bs��v9�M�JӴ|��[�a��nC�jT/�������f��7�Ð���ِy[R�a��d���p��ѱ�掙�I$~4�۴�l���V�����^-�Ln�����'NA�L�4iSc	x�ПmYm�ص���&+���j���q��d�	6cL�	�	V9�F��'ʩ��Mi��ސf�����n���ѐ	m{�V�KA�r.������I;�����zxD�h�l9��쫐s��P��ĴQ֥:9m��m�iMH6h�,ܯ�܄M�E��|h������C��Rӭ
�)vw3�ÊZX�
�D�d�5���I#"�6eCPaF��;����4�"�#�C�|hG/��9\�v�BY	�s�ib*��w�Bq;��>HcI��I0����:�W���d*_�^���)�����{�� ��D9c�e~��fP��-�"혎�O��d�<��A	��<<�
�|R�c|�C�\�I�9��i�� U�	�{<C�d���=��%m��z6�;&3��d�P��og���=��+�6���bƒ@JmI�k�����b\���L�&���L��ldM��Љ�t!1�_���� 9s�0��D��^�}�	9b���'��C����.�掞�);v�Ģ>���K૽�Z>W�;�#8|z,�M�$�NL���	�vy�cXq��i�F	܇���v�*O$A��g�C�	�g�S�O�>�~���pP�z-���!C�ѵE]3*����Ih��^��M.鐐�l���^��y����l�.c�W�^��ui�<��۬���Mb˞w����4���z};��r��I1v����!m�� XkD��z�A�~�w�صٿ~^����V;�<E�YZZW��)���h�Ōςf��/�;��BY(c��䞇�b����M3��.��wH��t>��r_6��'��da�U��|�[�yly_�P�S~���9d^g�6�IM�������Sive(��5�ﶷl�����;Y DZj�0�'��~<�U3�c[����g�6���g��J�i�;و�ۻa�`�4�񥱏.�����yBjvz��V�j#�)�_v/�l�:��}u���mҡ@a���O/���z>޻�����p����~f��Vn[�B����e�yA	�L�-}�Ki��P���3��R�s���ݜ��:�[�P�]�hp!0����2J͟A-��6#Bet\������yyI�}��(����!c/�,������!B�6�u�uxkD^k|��4������^j��`�f���K\w�O���֝�ٟ�o�x�;�Q�������|2��ye�>�evn��9O�����k�~s<��/^�m:��3��fn<0�P3� ���_��G�I�VM�Մ�e������&!�ې?]�q��)�1��$�[S ��=6/	X�N?�g������v�����z��eyezJ������ࢯ�~�'+F�n����_��n�8�`��)D�w����]�6�s�FϬ��#��Ҙ+ѝ�E:؂,��u/��U-`1�R߫&�zJ�Ѧ�9�l��=�LzT7��ڡ�`R������Ә̑��ç��(Q$�����
_�Rӭ���3:Q� �0f2E�x8��m+��X�O��}M���&Hk����R�=�]�%�l�K��G�//��F=�ܽ�=���V��~ �Մ��`P1��)���}c9%�����G'nˋ�%/O���ۣ%��ٚy����_��a.��T�q��+e�����c,��ˁC��0�͚Mp�����Y��u���}8��R�-{���Θ=f;�;STL�
)�n�+��9�>�G�,����+��${��
de�L�)�P!m-
)θ����Y[�a������e������).�ެ��o)@�e�P*�)O���vS�u�O3�J��7�C ֧��q`{������1��	xO�x�{��{�T~I8���}��8E�0�c"˳eV�5^*��ċ�8�K�C�����j'�&o�v�:V���e��&�)�zp��z�D���zZ��(��?O��}V����]Y�j�]kĴ���d}r��/��a�X�C�y�N���3�ՂIA�ӂY���t���@<Uhp������Y�[*���6��E%Ă�F;���y�k/|c
�o�a^��i��_�*8��7sa������ũǺ�����K^]�=�[��.�?��Jm�]+��cy�Y�: ̣I��u5�H��%��ü~��OHk@�yde�u�R<x\'ݚ�O'�ս)�9Ԃ��v��\c���@s��[�Ī^�KO#�!`s�8�v�f�������k%xL5dy��������=Ff��
.�^I�2[z�ۂ��Ca��.�~��<%`\hC8�gM!=<�	K��)@e&��x�jy���W�Z>��w���^h��)ќ�/)f���b]���Lk�,bt5r��9mB�ZF�A�q�Ď����~߄�z�B�^�UL�3�NA�(a��hdXE+5��>��xڇ����A최�[��nQ�/c�,��1z����I�5�4ݱcÉ�ː\���
Z����gx�b>�^� ����<M��8ϒR��_Bf����f���@���n.�k�w�$ʦ:,��Bx�p��v����&���͂y���]���C����te�^F�.k7*����<�]�йώ)r���/����� r�)+�m��e�ttc�K+j�I~y_����� �����(��,��!�b��c�����7���'�NJ�aj�FR�>&�i0�u��4f�D�㫦#���|������yt��dE�� �qx:"�S�>���!k����^Xp32��I�3/��5����]V���-�=��g;`��NwF�!�nZ��&��yyήy�[��i`c�=1��=�x�DW�{�1Ǉ��@<��6�x����a'�\~I�{��z ��g�_J�Wh��3� ���Ѝ�h��zՔ����,�{NxLB(�{���rOQכԆ�(�vz������������]��>��o��1��G�^г>�~�,��G��G��AΞ�/�����W�)gyڗ#?o2�*�G�dI���iƐ�A�Z��O�bbp������C�l��0#�c�֖R��1a!k�{ȨV��3�b�w<��f�S��W6
���7~���e%��
���	<����(�\TX�0�R�!��S��ă����h�I�ƳQ{�[��gX�z��w�%Z;PQa�����?���|=_z|��}����������a-!FV��Ɍ�e���ѥ�3��~�4�o=yKN`2W � Ӂ���t�g��^L�U���5W{�h�h�<���$m�D�Tj�#׈��ۄVNȺ�8!�B6;x�R��]�9���r��4�w��	;|����{���{<8KH���k�#I/O�/X�n������c�<k����g	�a��F�Υ�\�8�1�7�I�{B�����T��4�=w�]���]�;�����c�1���py�o��Ɔ]�b'9�S���j�d�#�����"���s�Ou2e��+=5m�{^-�JvB_�S��u���CY'�wa�z~wύ����]��ڴRZ�6�D�E��:��L��c�4�t0P�0O�*f�4k6K�%�=�03�4pá��!�c��}O@aB��1IPy���JO����	1K<�g���s���\����٣�$���29?��ס�W':^{Q0���w�z�Y�ג��jM���=6^OQ^{=by�ǣ��L�^���!�p?�G����ychc���&[���Ӱ/]�i�����AC��<&z���~V�R���l�׎�l=�./nX�*�fZ�Χj���1ᇦ��d%)�)��/�B)jg�q�C:�H"��v�������SR���8�%ffܞ><'�Z;���I���w���B��ӫ�G��y��}�����C�%��,6a�_�k��.��z}�|X������g���"�\����[t�?�]MQI�Y�<� ���t���$� m��T;E�ðM�l��� ���:��"Y�6�u�qճPN㓥F93w���sV͝�s=���.�B�f����	�B�/&��K|��!YȕT�w`)[��LÄ��:v,��IT�ƥ+�N:-��)��@������̚Ⲽj�������=�ʂ�m�(DqᐑD�5�G�W������X�5xB?\ǒ���O�y
�K�r��� ��V~I��?׋�9��A���h���ۈ��;lE�{�������^��#�
g�"�͂/'�E"MV�6cQ�/����t{6�>i)1�K�v�m�I~�zRN-�F��6��U JD��*�[�y���a�C�f$�Sy����xH��'o ��(�YY��7��
��+�+��\OY��`��מ�^%F��<���H%�g���|O,�����^��.f��5S�|�y�()[�͞����$�Ƕx�4��:�����KTR�Ы�I�i�FP��!�w;9{�,l6�t�rH�%�͢{ݸ������#���>�5�t*�3��?�v�gaZ���
H���B/�H�5�o���T�z(HL!qw�=}����┍7pu��������5����:>��� Fe׸�����u��K�Ɵ�x�M#���]=�?�Z�T�Q���g��׍�E�����&�y�pFڰP��졆�+�˴��޶�gC�L��a�����v�	]����>���^��m=�Rj�QG�ʲ�@��4��ҮVy��$M���m>�Hн|��X棕z���Y5i��W��"W��D����>�5�ǩ�ք����p9��y+q�wcI�B܍�-ʙ�O��{����KM�z�	R�J5fr.��{s6��0�υ�����ݘ�ݰi/�U{�g���.4"����_�C���,��g�������ғ���
��\���၆=����X	yH��\2��oOAx�҄�Շ������	M2�D�A�ܛ���b�	X,�<�94a��x�lb`�IBeoe��W��`Ss���o�`X�#**k����"-��;�+ ��|7?wT6�]��B��1�μ�°�ט~,�S�J�Qkg� ���m����A��`�=i?:j`?�3����<��xo5�7~y��兀^H{}�r0O2笴-���^����^�EX'�ю2j�`|�\?�4*�����X���qv�U�D���s�?ʣ~�s㛟�_�y�o���6<�݄�L_��~`��[K&hb��,PX��6���2�0h�\�4@�kX.��Ҡ�'��C|�wKh��w�<�`���������х�^R��\������'��]�]I��l�2�d�v*}�zx3�9�,�q�ݣ)����8��� �,o��Bۛ	x�ҫ֋�ٻ����xľ��.�Y4헛�r�P�Z�9.˒�V�Z��4ߢ��e��.۔��x+���n=xBA�AdШ�?�sX;�����払F��s@�VԅJ�뺵��Mgۦ��؊$�n6y&!�d���YS�N�.��$��<ff!res^%e�	Wo�qJ=X��� ��G�R��;��Q�y��Y��Փ�ඕ���hS�����C����g�)�/>��������*&�O�{9o�g���y.�of90�ܘ�~y*[�w�t���'�Le7q:mN�,䪴Rd�gc��Ε���}:el�!���o2ݪ�W��zf�c���3Gq��$��i���Y�Єc锁ZC�8PNM5��P*d^��6�XFj�yM��������{��X�%�m�\��ip/�a���R%�Ʌ�Tk�%+�3����6|�����m�,�k��O��������o����8�߶����sr�Iyu��M[H[�=�|b������qU����qv����K����`�SvH�5��;�����N9b�A�����݇p�:&�b�橓�<����^�w��m^9	i�[>��Ynq��l�7�Џ=�	ϒ2���	Z9�%$N�~Fu^�5a��J¨d럞+��6��7/�{��R�����`��/�>��T���[�F�7�3r�=G�����8��\�R<Zx�T�6	�VO���c�[=�#�Y !�$��}�-�}��c���1,�Z�o�b���l���−Ǐx5�U��J�	 �:��#ג�Ə�0iH}�M�K����`�Qx�6�"�Ҵ�t��JL�&O�֮��?�Xx��L�v1J�2j���d��S���(<���<%r���~)O�!�9��
��Y@�������`�=5�^�۱w13َT~����1͖�c��i����<�XQ�z��0�~�k0L35�-=�}�(p��樊EB�H��Vb��t�[k�'�dWJ�܋�>��^l�Ճї6�����Iq&󯷘�w'&-(
�m�r,�6$�Y�d=�@�|P���a�Jb�H\jE�y��g��>ioR<0�)��������0��?V���WM��3���s���1}����S��[�JJ�T&��b��yʣ�޵�����þ9���)9��=�x�N,hu!��\=�!�@^�h�y��ϕR�gm�2Ek��+���i��5X�a��4�֌vޓ�q��JAME"�ڄ�ӌ �ѓ���]�r>�X�+��fe�n!�Mr�iP"2>��'̃gխ��(�<岗<Ġ�<,����6�<��=!Tb�ڠ-����2ypym�Cg����=A���w��yi�x���_���wt�!���3 �	<�
Q4
�R;=�t�|�k>ˋ�e����o��1m�R��%y]}m,��=)^�1q>�x�1@�v)����,C������y-	�e��u��
huhP��/2ݪyG���hTk���)@���mh�1>��L��to�v�ů���y	h��H�_�qW[�kq6o�R%ӎ������4N�z�0��}��niaZ(8$qǔ�RDT�PXK���^����[dx}n[�x낌k�2�{xM#5Ԇ�Ą�L�s�x�r��뛓@��?쨸,_��4�3zy� ���Z>V'�)қ7����k�G^�fjB�Wi���ST,O�co.�
��P'n�m��|��y	���m �@'ߑx|������$<� �s꫕�ѧ�:z��õ��ﷺ�+y�Y�v�d�ng��҂�:�v�̓t��� ��*�<;`�n�磜;�?��ۭ���+]n2����iW\�w�m�������vR
������a���!B�	({��<�Z*=��{,/	�v�-��N�)+�R}y��^3A5�z��86�����/��W7O0q[ysҔi��*^ov�m.!h�L#�}i�-�Sr%>��y��-�w�τ�����S�xe�~۵��O^��c-ݚ����؀d�W�|�,��W>��y�������ާy�~2G�F�+�i��t��N�B��5�49�K�+�z�C�C�k	����C�=��K��6K�+�ƈ�@)?���f�K�+�O�9/I6�PX�0���h�}�G^G�k�J�̳+l;fV*�6O(r�=��
0�jDO��5\(G������嵹�J}<���f�a���1#q�|����'�͔��r�b��m���MQ��,���9y��FԵZF$,|ߏ� ٢�����n5�N�*�O�Y$b L�$Z�i�}�C��z%v��c/���c,�^C}���*��%$��Q��:����/E�{(0P��!8ر]l�bΨ��=5�x|�kRv��h���=��6�Z�u����+<�΂����i�<O��xb��k��ݽ;Θ*(�.�b�CX.Z�Iڧ�悙O�29c'��\��J�hRpÒ>�w��ք�f�}2�N�&��vSw��5
�[�����4e��&y؎���۰j�B@����J�N�I7Ttaߧ�ue> �%ܐy�X�P���)B��;5%�l˲~��J�bI�\�}5%�V�ʴ��Lb��}NYī%춉������/y��h�ex���*����K3 .
������QV�x�aIa�}\���7�d���ȧyUe��AP�J��ZS����WM*{H� $9�L���c�������ˈL�$�%�1J��N-!rV�|*�r~�q�:;��zh��	�K���:�c&1�)B�CY�~i�r==��]��3��,���J��{u�T(���+��J���N���:��RH��%a�ӆ7'a�(�xQ�{tb����	욢(��S�(�n�瑮%`P�/��{>�����ܸ-�\<�\�ǞQ 9�iW�!z|�~*��w�_ʳqs'�P%��]�?�h��"�}���KM����mg�c4񾑓�[#���(]�k�<�3 �����_�aK9y��m��5����y�����b����#-�L%!X0��%4��H���~{�ՔG��^�J�)�U���o+	m�����tM����D���l��g��|X��=/_Ȟ`��]���{̣.^���;��u���V~	���6�<İ���Ǖ~��|E�ɷj)��y{�E�6,r%N�J�6��`�Z������o�/���(zC��������0Πw�'4�Z8�I+����m�/���j���&`$r)��,"	{��_M�z��r�7�e��_�s�/k4�A�Ճ]&9������`b�y��S��{B�C��B.׻�=�g!�
�D7�ߏ�'�Z�Ay&,�������>�w��q��ۥ��_[;V�䦟y/R����	2;�+����d�+����t{�;W���uf�Th�u��cagc#7!�p��s!�]�ّ��wJ��v�ϵ�gI��	�ب ���6ͳ*���&u�Bt�y�zM�ɯ%oA��3��uY���S��v��q�5�8f��U-����=�<�x-M�N�Z�Z���<�{��C�I�&a�q�џY�ž��GL�z��:0m$�`�x�����S�߲~c׬nbS�B]FLRªmm��v�m�ѬIv\���2m��;���cm�\"Q� �A�kG��C�[���?سVW�#��<�n����B�����=�}km�|��}c��� d�!�_��i�y�m��=n�IyY<�FyD�#�=u�h�}8�υ6���~S���4iO��x��x����{�r֭��z�����يP?~��F�Ջ�}��1_3�|7������AO�?���a�e��}��������a���xM�v*��)9HS���1D�?�pɸ��~��D��(0Ռ�<t�����{��`�̈�9'�1x�����y� �����F#@�>oö���&΃���bIZ�,���3���ԫ������y��V��\.��)]L6�������(���S��<�r����h���H���t/#w]��c6~~��4�(@��Ih�%���C�#�:}�K�[���H�1{9"{A���m�v�����+F�>b��}s)���nM�ٌW�'g]��B�C��֩tϻl�"��P@����\C�^����FL�,���2ͳ��r�>��gm��W/D�|�GZ1�K���Ք���\/��8��B�´�>+M�p<�xt��Kt`^f�͊C�.��=�ym�gj����eZ�����5����`'��˹��7π�o��Y�C-EuB�5I� 4i��z���!rn�d2 �o頁kȯa�<�����8m��i�M�-_�
[����@�|xPc*	��o~o�������i&�Sx�Ў�6�|����W&ҽ��K}Ă�$<�)x/�#ulWɣ�i��+��|���̦ƷL� )���qY�n��\�R=��Z2�R���}��N��t�]��4,<�$���C�R��8�D{���t�H?�qcIs&M�G�I��a7RWΖ���jC�i+�C�D'�M��F����0	kHO���ufȉ�s���%�V�̔�li���u���|��Zb�p��7(Q�rL^�=&�<��M�1F
��Ѷ$�ٴ��)�2�G{7��D���w�,o��h`��ă��U<?x�cz�%ŀ���R�,��J�^ݙ����ﳒ��,���F�g�'�\�ؤ�j�o��W����%VX�D	�3�a
����C6nȸ�3���c����:��2Bx�rg�;\�:�" %��y����s���"��eƶ�-D��������`�p������C=5�RClXO ��:�҃�FA���KHޫ������L�]�������l�%�����>���pF`�x�fO�`[ju-���X�3��ߝi�uD�\�(k����S<�8?桢{.�����7a�>��Ε#��f��O����΢\߇
�7
�S�˴�-����/ߊ���QA^��E�f�
�Y�Q̼�}�cF�b�eخWaՉ���m{5��uqd��t�JP�Y���nB�2�0s�2+`�yY��p��g~~i/�����7Xg������##�{���^b�'	�²JH�d���{��X���vl��E�MΗ]�6f<���)	l��n:c�xueO|���{�G����������˓��x��M̓K���A�k��<�Z�~�d�K,���}?����s	��i�1���gg������bm�⎩Yh�M�5~}1����'���vJ��;B�?����]�[]����i`vܠ6��̮��t�9�k���ޘ<a�=�m.�GFVs)��J�$��,c(/�;>�Rn��� �@�lBa���d���`�wK߹_����_C�%E���us�DSԄ�iM��3��Mt��"}QiX�ެ�ğ5�Z^N��4����6�z�GW|��� �~��ͱw�f6��5�m�\%[~�%�i��c��'% ��9ߒ��M�.<�Rӭ	�˫����v+6������k�>6^�B׈�eB��i���a��@M@�C��T
ʟL@����tJ �~���<(`�Ą`r�\�@��9l�ߴxK��	�C�Ԓ�ٓ�녿�C!r�,�� �:Ibs���ZS �}���%l�$��0�����X e�;o�ܴg�H��Bl'�X��#�Xp�!&|�:rl��aB��Q	M ^��3^Y�<�bc���!�xB�{@���؏�\���F��ntZmΒ�XI�����z9�JB,��@n�&/�>P�C�i����|p�gw��>���y�1��~��Hϼ�j�E�I�Eޙh�h8�͟��]���D�U��P`�2~Iw0i��aLj&�0YbV�Ɣ�M��ī��vp0�k����ѡ0����P�Ԅ0��28�Pf��J���%����yF?��-\����d��J�e$Y�ǫ��c�:��k;�Yo��q,�������E	,T�C��<k�y��x0�x��̢�c�����k��l��(P���1b��`�=<B�x�]?����� ���n�y�8�2��iU��bm��kb�oR6IB��q-杖�d�f7�g�$�w>"
N�N��s��3�p�EK0��3=�@)	�D���
���7Z2�NU�S*Ǆ��<���3%���mp�l�5;lIA�e�9O�^W��öa*ё�h�����N�N�6���X����'Ao������c7t�{v����l4���@�%���r��;v[Y�L;�ͪ!��V�i�I�p���0cz��%kx�2	�׿��&-�g��E���ދ��γ�1k,��y�[K��<%?��ҵ���K�Fy�Z��2ZB�5ŀ�q��u(չ$ �:�O��dI������^�O��uif�j�����k� ��o�_>r�Ԇ��c��k��J��{�4~<a�).�S�9���kf��ֳ<K<6��R>y��Q����G��N�����D�A!�v�ZJ+���3"��I�$���J�`~��)���
���o��������LXF��F-yhۏ��@6�˂�8u�z��%��|�	?�	Q���gj�'�P�3<a���\7n�ոM�x�J�T�wI,���5a��ͧ�c���e�p>���p�M^�%��J嗒�7d���9�QNϒ5����"a�}��*#�s�,��G���Ot��Ї��d��c�a�I6Ƈ�u7�{M3�@�wzŘ�4���;��
N��96��@�g���^5%��y����[�=�0��^#�q|ף9>[ʯ��K�i��ҫ��XYǄbi1��(���x)����$|
�����Jm���,̏���*����2R��7� �<k�{+��M�,��9��.�w��׋M�wr�H��>����7��m�z�nD�x��#�Ϻ�c_ĴŹ���>oc�ƴ�ARZ?�����o�^��Xx1c{e�@2&b%���8��5v�u�>���/�qD��_�X����7���7�[=1j椐����l��gz[_))��RG�W����J�Ɨ\gF�~dD�����OX���hJ���!�9q9�NB3�g�w����;�I b�v���Q6��t�Nw�����݇�i�<D~�}�9[C~��RR�!��s.�bā������l�Z)��o��G��ʜ��#���y�sT��I��%{�c��-+)De5���ba��g�(|���@?n�*	j,]H���w�����٭$��:!�NE����ѮV<��}�=[R�5��:H�!�&�,����]=����G�mC��57����Wj���FE���]��&�7�ݰiӸ�m7"�Ճ��cc6�j7�?���ذWaq>N$������^�=5j�gF��
���]H�ΰk?��H��F��\�+	�6j��wa����n�	4χ�Ãpvv֍���r"�0*�,��W�2��g|O�x~Έ^�q���3����n7L�BP�)���o��}�M�.S�R��o�]�t7ee��+֕)�q�uX�b����y���ny{�Q����=��eH�c�:b�KB���7s�m�4�x1V<^c��s�hB���9D$�h�ڻ�F�����3	�7,l;�oo30�gmϿ�̿�:��u3T�&�Vd�W^\.Ȫ�$�G�o�����v��j�����?X��|?Z���#��QN$:��O����~�g�QN��Y8[���g�ec-Fv����K��b$�Eh�6l�U�jQF��,5r;ʬ��X�㣬���ۉ���� �{H��l㝋���QAvd�%��x�eS0�4�$�X��Ǣ� �܈bG�� ��1����U>��:��[e�ޑ�X�c�B�wJ�1��V�	Koᓑ%^�P4#D����>N���(
褐�{��P�J)�-p~��󀍫�]��dP!{30ۑ�NK���hp����7��g=0���ʱ�XW�x�eq{=���~����K(�
�4��ȦMX�i���cVb�ç�՝�Pr�t{��6��]%�T��}Q��,`Ԯ��(Uv9��4�U�%D�-��}�	�9Q"���6�<|�ڴ�[:M|d'T>$��X2o������1��gj�þ3R5AlqXx���_��32�ou�gl�B�HD��>�OI��uϋ�hMy�L���S�6轺N����uΫ��̱���H����F�^�?o��W=�{]�u�V�<F�Y~��x��=p��=_�-w�7ٳ�����|�<�?'�a������*�C
�K��g�KM�zF�!6L�bO�n9�u6���ҡ -����N�<�pes�W���Zy5T]��h����{7?�#0̛�%Ә��m-	��d�y��%	�M9��w�:�Ь)3��m�+	pU��\�Z���b��s�'tJ��{<��W/ί��\�7C(�.�� �0�M��
 �9����g�
}V��&?�Ms8�]��&����7�n�`t��.�K�]�rW��񺜞%��ρA��b��{D��?YgH��Vl�ًd�]��,A�<z�"0�
�#��C��a���ޏu,٫�p�6H��c]uɣ%)	gc!��Q̈́��������{��<��B��=�kǄ��������RV��P��IO0z�b�u������
��B�pM�����s�Ϟ���y�xJgـA?�F$�ք�c�t��0D��?(�����Sm�.���
�gE��r���~3:�fz/6���\Iʼ4h'�/�R\d�ȋ�vd�?�`�u��l��������h�AF}HB�x)Ό��SPf��lB)��R��}Rr��������ϳЩ��$0�c��~O��s�..ӫ�'�8/�,�Jyym)m�{���h�=���|���w8f=�2�����������y<��=�R+��Lk��u���b��M�#������D�M��w�0E�ɀvA���q�q	��y��v�;��5�D�Ő��d�!��'���c���fYS�M	� Xer�;pc؎���e>�+�L5��P�m��^��!k��9F�,(<�Ech�(lQP�:�����a�Nat}2�ۙ�-�1���PꞐ>�H�l�^����g�U+�S�UIu�PM�rJe��y
��6N�{������+����gP!	A��/?5ӳ�_�+c7�/�^ �  m���<���MM��#=X�u�tX�
��t���E�6<��|��V��w�
RA�\��)����=B4Y#K�i!4db��w�ZN��?�^�0�ߟ5�����if�9h�y�����NueRC�ѡk	-�]�ӧ�6{��^B��\-o�7��	cM�y<��=EQ��1�T�=�8����}�>/2�f^��������>F�z��b ���x���d��&����~�22�k����#�m���Ź�'��jZMP�r/Fh��O����t�e%zS���K�U.��*i`w֫MX	2�x�z�G�~x>t�E:�F5�H��.t���}��a�?_�S��xm�j�P��2-DI�kI���K0��H�Q˹�c�7�����'1ѓe���s���~|��|�+�<��N��.��f��X�cIw���)lC�Ӝ�-���E~��>�$({��aĨ���^�O�Q��U[�wU��E��y�y�����v����ރ<h}it�L�GP!�(ƾ�� ��d�@��{��:I2�~3OY�}l�%���B���o%��>��6�z�]����n}'\����P�m�!u��Y�����0���Y�S7��Ժ�rx���N���Hrɮ��_f�^�>����y�:�6�H�������U�ㇱC�0���V7_L������u`L�>$�N\2iMۣ��TB8؆t�B�>o	��T�ӵ����^ۗ��G���9
���rQ�x�*)�\�cȓ7Fq��������Zº�l�M<p�i��7F�S{�g��MSX?�D2o�����uel�D�6�"�/�֛aa=�B�<x��{W�Y8�Ϫ�6���8N��V�����O6�.��qj�8� Ȋ��2�z�}����;#�N;�bة��(���N���!�9wύNV�w!f_X�,5�h=�6���|���{���iE��a�C"ر��䡊c�����2ǁU˳Ĥ�2��}����A`׽���y�h�O)oV���s�:��������
(��:�+)���z`�@a�)�R��OQ8/�`�ˌ���/��x�gW�����|�K4�ѫ���5�D�u�8�N-چ|���	�j�\�W:��u�ÂCta+G���чE���+�(�B��t�.�i{�GSnI�m�������CW`��w��q�54�Mل�:��! F(���66�2���fÍ�� >�]H%�ϔ8�+	|���|�]��ZY��ҶP�����_~��&
CT(^~\6"gK�S��r /O��kI�`9ǔ
+n.���{ϕ@�1%<)�B�ql۳g�j�%���v��	��� ~�Mޙ���]�!��7�]�w�Z=nl�i䘘�#��$�D�Ӥ.OsV!ѤI���*�ͪ�l�1=d/Oy[Q�0�
�4��]�8e!LQ9�ZN	�z��RI��@��28����'(MiԄ��BB]����<dUf�A\jq~�C�^[�s�ԏ�.ׇ�!���Q�#�?&Լ�X�rYh3��>��q���%(���X�#���qV�3���Koܖƞ��5���8$�C�����lE���c������{=)p7�Ԭ�����m� f��l�pև
��t�~��v[ �1��|=w�4,B��G���Z��a6t@��.c�Cj�/��C	�<���c><�f�t���R�򮋠�',Jy3M��2��	$��M��\RX�� ��^�]����<:p���P<>���J~�\�c���c��9x4D�~��e�񈗎)_L��w�م��M��P	a=(�,3�;"�Ж�G䌪m3��?DQ6%)��֯�#�Vۘ����X�C�S4M��H�NN�Ħ&qx������Zv��Y����bÐ�.~�S����1!Ϩ��Y��E��=az����NA ��7NA��\I���偃�tp���Je�C��u`Qxk����K4�<��p�֞ETX*��`���ői��A����0i��아���)����v��R��o��Z���Oޜ%!J��^���A���t<Zmj:�a�n�*�(�ؖ���w���y�R�ɾ�!�2���۫�˦��e d#D�S,�l�o"�B���M.�ˊ-�v��ځ�I�S�U;^�O7x��A=�l�=%PCr2%<FG�~���P/���ն��3�.Oy�q�=af�#R��B��ӣ���,8�,Aj%��'@�rY���ҙ	|���r'��S�+��s��]g_~�k����:�8Tj���) ��iL��zoո��+[�[o�*w��A�:�u�Vv��cuv^��M���9�pw�tkB�J�>�;۳��r.�n�s#Q9��~D��/B�������Q��>>P�ə�z^��Fa~G5c/����a$Υ��l�����p%�d�ԏ����  ��IDAT���}xL��ӥQk�{i�E��Ş�[�UK����A�voF7�����6#Ĺ|J��=�O����2�
P���a�Q�g�\�ga��D���������
��W��)���
�}�9�'���|���E8Z�^Tz� yy���T��!����b���v6���7\�`Oރ�)O�\�������x���]]�YĮ���i��b�	��˰�G)5ʧ��K�J�Ϭ4��X��>��Ja��J�����Q�t�8Z]�}*ﻻ�]����V�`u+��j}.�!Eg�s�����Q�uM�Z�:܏��~�}���8^l��3r����#���Zj��gbTa��V��0a�Z����t�X�K;r�"^�W�����"/�e|����< �r*	~,��S��(t�:*�Z>($ya���ނ��?�~��p���2�՝ֻ�=7Hy���i�3�®q�3
3o�"u�������ǖ<i�����i�P6#mk��Q�A.��w��{��������&�YYqYX�x3�c������t6���͖fd~��S��̊���7�n�es���&%�|}����}C�43U����A����������Q����ӗk����u��3+=aRz<�F?l{�L�$�جČ�4���|�P���/6Y�_���`f���b�[=� y=�����B߿_����ݻ��,�Ƒ�V���#n/~X�6��N:Kʉ�,�~,��g[g�_R��g�W=��&�``���װ��֌�k���-�#-��p�������錄ɿ�J~��4I'��<�ۼi+T H��E&�O"1E��$|tyyn2ݪ�&��t���9 ��{B�=,Z��N@.ii0�t�;5/Ɯ�t�=5E�ĒK�R����D�y�V�[�KmB�=���#�+���2=�fHK��⾕d��E���T~�p�k�<�T,y��[�ĺ�@)�����`�\�ͳL��u��S�F[��w�v��<ʈ�6K@Z���T��ۏ�{��ʳ���>���6ݲ�[���L��a�j 14�؜�� 2�1��x�Ƥ�ر,T�˪���E�t�LZ�'^�x׃j�>i��3ɜ2���y�Nβk!�����o�b�T��_{�6X=AT˓N�#r�X��e��Q?�[�	Z~��G�޽{�T���|F��v|5:b{�~H{F�aP!�}���GӒ��~b@A���3��ݣImLԐ6*�Zbz{���{\�wM�|\;���^o-B�֛����a��ں['o�W;��N�c[M_�fi¶�C�/�줎g������ҭ#}�[�
��>I��]j�ٌ>����v{b����OU�>[N��3��Fk(\=��1fi����)}?}QI�p�<p��r�
v�]�����b������px��_����x2�����/�� �}��-�ͬ��q�'lA�򔩸�C��� J4��T��'��S&^�2�5>�wk�g{�b�f^�����Yn�:�
|T�J�����L�MeOc�7����Y1�Q��?��M��_F��w04?���ڐ5���N�Q�/��X��(Dχ�J�,�"��Jh�ʺn0��֙��$^D��=�`�� (�����K(�{����\wdf��G��7�`��՞��:ۢ�ԏ}�c�W~�W»������GѾ�GL=b���4��A���Y����2�,8�3�	��G�[�����7�!����
�-�z����k�ݸ����ü��keq~<���Xj��S0܎�����J¸�;�4>�M��<O:�	y'���t��oT�!EwU+��ӹ�!��:�̔
b�P3u��t��K;t<5FR���L	����|̦o��ɷ5���<׫�Rp���s�;���,��=��ױ�p�5;=h���ɼ�P��+y�Xµ���o|c����𖷼EQ����nn}�	(��˵wJ�����H��b1���O������[�~��~,����'�¬�~(���j���i�4`�ص�~żk�֫#*��1������k;>����&t�|O��6y��zx ��]Km�'�a}��Zݯ�Wuhq��|I�&���e� ����f��&��f"���߾h�,@�'y���Հms4���ߨ� ���!)�&q��l��c��g�"�O�g_n����<�LiXbc��0�w��N��<(�,�9*UVp60������/	U���;��FлrA��T���_�����9�~����#�<�e�o[�~6~�A��ce���A��G>R��)�}�6��K��K��������2LQ�����m4d����v�b��fvµ�V�^���̧�R�	�7�Y"���@�/x��ļk��c��,X�uX����M��(_������[�'��\�<���&o
�颊��w�Jv�&���Yp�b�E��+m�4X����4�}�����hNDz��PF�me�4�6����Ǿ�G�>g���(�N!����?
G~��J-OoM���h��zu�:r<�Pб$y�0�(��&�m��������~��>���oV�/�e/{Y���?�BC��pf_�:�Cp��<{*j11�l����SO�W��U�c`�B�4;�:1Ͱ<���B�!	g���^LT4�~���ߵD�/�1�>6��r����
�\ƫ% ��mv�l@��+rʛ}h>m)Ә�z���s:�t��t�a��C\���]����x�4c��J�tЌ�;f��oTk��j��NΫ�a��4�I�������1�e��!����و�;���ٻ��J��Zb3�'l������{,<��s* MhJ�ɽ/��/	��˿�����|�^�ԧ>���CF�� ,�+��У|}צ�Ƌ�uO�zVLM��c����������i����L;�f�,�Y�����yz�K�8��pP6��fB&<p�%n^[�2/⬔�JM����9#�q5�Q��01��o�~�d���3�_�6оv��eS���!]�����i���M��2޴d��9�:=c��lR����^�|-�a=�`��pk�ѳ	}�=O���X�7
�R=k�ǙBi�r���R{����O�?��?���'�;�����<|�W~�
��~��᫿��ß���{�������1���W�گ���׽n�]�����[�����֥�vĢ(1��moS���w�>��0��G:��X��֣um6s,a6��fw�T�	���y���+E���7��
��K8�1�ye�M?��̮M�ĤL�7�B;���w���M�>ؘ	a6�5K��M�[��o[�����foӛ죚${�)W���T3Jj�i��p�X����4�-:v����(�f��yPX!����Z�0��a/Ms��1��	^OI�[-q=P	L('$!Cy��z� �������Ї���|Mx�{�~�~*���g��G?����Y����������!#��� ��K�{J�������(l䞭�X^����U)	������)��ңmm��I��P�� �R?1�] �p�k�sYlr���.�����Qx"��s9@�T�C/B[�f�`�y���z�n����d��iJhW��P��3��ciH;�%z�����m�;5��!*sg�ڰ���Z\)+��'!6ђPB�L����ǐ3��F�'����w�Ց��%�+��ays~��`��^b<o��^��� d1�|��}_��o���׼&|�����E��o���fQ��mߦ�⛾��}��W���j��E}X�����W��jB�xWڼQ�	O���%�;Җ?��??�C?�$�rM�G�N%���3��u���)_�g�)v��;ݼ��>��}(�1�_m�rٳxN-��@e��,�S�t���e�لyqZ?!	�صy�g7���]ȕa�-x�M�[��#Ahq���`㒔��h��4�}�_��t�{Hv�!��W����-�!��+7-��8�����P�A�B�����<8?OP"2�Ab�-vw�Lo!��5�RS~%�"nG)y�����s�+�b�!*�S���w���b���o�F5�����������Pa/�Z���2 -��-�z�TW�<�\e���O)K�&ο����)[_`�ey`���Q(��b��;>3�{��3�yt+����J�W~���T҂�RP�%P٨�ˑ��4��O�s��v�ʌ.�Q���('k�y��d�H��i����C���{�Q�-T(7$ژɅ�|)��F'S���΃"�>���'�;
�i=:x�f���{�<K?}��z�F�yFQ��X����b{xIPab!$�`����œ�Н�r~��TO�����j3�@k�!|I2#�����:�%e,	��ٮy}g��|���˩������>�ɟ���V��{���wl0�l��$�٣�G[O�r[�v��v{eK%@�`�x
����"�za�p�"  M�<�f�{8�2��Cv�	�or$�U��i�O��c��2�3g���$@�z�M�[��ͽ�C�\���}dO�U?��u�����K��՗�5�I�>��]N�Qiԏ�WO�xz�\�!�FR_&�܏�JN��.t�f|�B]���+�%7�����gMx�y>l�GCs>�����i�d��ʮy6�%�馅��g���3؂�5['���P�ZY�DjúX^�'�s��%Y3H�;��ʷ���ei0Z�����|`�a	��C�!��4_t��|n�T���������*X�kGf vX��g�����J�]�>4g�k"����4#����������u!A��k�����n����
y��I�3@��B0�u�'��	�Wha}�B��������LC�|$_Z�\�S�~l
�w�?QY����ʷ�X������ߛL<
y/f	��L��9�Ġ��(���B�݆�z5ʥMx����+�^��3�K�߅+)�gQ��UKq^��l��?N0�c�X�u3���A��$P��G5���!<2�~v?��G�5�o�W�h�c�_9��W�}��a׎��QD���uҭ�a0�S�t`"�FJ��C
x�"�oM6��*��&�6�B�m�H����w㼇B�)�,D+�3��Cz��!�S��<����<��f���M`�g�	l���>����V1����k1o8O�+��*�0�O�,�2�����>��O�7��M�g~�gTQaB��<���R;pO� ,���|<>(�B�V�<��7G:cY��Ʈ�561�Y��s^>����{����$����s~ͤ8Z��!+B��ŠQ�aT�/2���;�f��i����������H�[�����\BFa
�����{Atm7M{��M&�}���"�ɠq/TH�;%���F�3!�=��M?����a��yJ���9Oxz���K�P��+�$�9OF_���uFd�pe3{�s����N�l#�a�=��Q-K���e�/�wv���]f*��X�&������-����^x�;���˾� �������J�R`{$YXhV�^<�R��~Kb?~o�p��;�u��J}�e��l���Mz�9�Și)�L1�<eȠ����$�RK��{��V	�M�u�G�}���X߮����3ě��e3M��ZX>FN�'�:3j#s�@��2K��AfFA$�e����,Xʈ����H��C��I���u;����wY ��<:����y3��
��ߡ�|���/�Z��5L�#�5���9���^BY5���u�S�仹���=[�Ǜ�W�/��Ȍ���{��
�Y{�y|^��F��V�d	�ʵ%{;�^Ya��.Kj��?�]f%������7�����KI�jޑ����ѝ��^^�`݄�|Vg� �r\�����5U��$ϛF�h�+���l��z�����bH)�Iq��!xoP�f�SR9� �P�7 -y���?eP��oF{ȔL�R^��:�еE��Q ��h�xB\�����׫_I���"+)[�{8{5G\N��~Mg��l� �f6�`]ДS����R "/э���7�<������kE��i��F�3����cVxI6�5�&�Y��D��S�$�N��|�x�j���K+��P/��ʥ�o$0جU.�����'��(�.gZ@��|��V�I,�Q�����1x ��A���KsAtP�^g���V�N���)��^CZ�.��>E������р��ϰRbE���"T��A��\.�<+�����1�nn����<��G�ZB��b_�P���l�T�$���� ]=��?��7{��x���ђgi&tY�X��7�v��Q؟^]Km���r�v/�ɮYͼ$�"&{P�֟d�'WM�{ڃDp=L�F�fY�J��B�2{l^�O�i��@ɦd�Z)��l�$�=!0!�S,����P:�?�6-�.�N�S�@�!�CD���]Mȳ`�D�4F��x�`ٞ�}�m^�k
����X.߮K���Пy�س�ZkñY*1t^ٻ���F*�I��MY��iI���7�9E�K�!]�O�
�=n�nlw�}�M7�`<%�e�ov�6x��
���1��]�L<��y樻l���4����Hv��yuQg���
�Zd�E�6y90�������V պ�� �@s�w(59rp�?!����	�[�w���oCrk�0���:�d�qvP3O�%�5E�]�� �	6i����� NU=�_|��gP藄$+�{es^�~��-�j� <�ּY�]�2��_���&�<�o	zƃP���''���r~LOU4!��6�Q1E������Ǹ<%�V�����U�g*�>/Ou��������-�ήq�c��)|��
Juc޴��G��_�k�~��S�y���ez��a�a�*]E.I{�a��X�l��^��D�U���s��U�za#���0�_���>ܹX��8&Dr��!{�hXe�F%���v�f/�[Y`iӆ�xv'� �y�r�찻a��ݞ¼Y�4����!s��$�͏(�}�-oT8�<���`و�JZ��1<E�mb�c�CA�XW��$������(E�s�J��)O�2�5XDf:b�{�@�嶛)��1_�{)ғM&V?�bA�v(;+�][��� *��'`M9`?���΋�-�x�y DۗA��a�e�Z�U'��ЛӉ s1Ew��X3"�<��K �mz��۬F��O�/�l5>#3�hb��=ǣm�nt��>�C�Ҡ�7�h7�a��t�Rb�����mG�|s�nM� �w/L�oM�\�׃'��i� �{ٶ�X��!�r���D;>TyZ�6Ԅ9��N>ԯv��:D�n�U;�����-��\�+�>�Jm:�>\�7�y��R	ɔh���¿��e%��������BR�S��~�ͥ�������<Zy4�zt���+ٛ9��	��3�԰\�$<D�+�\RKc��R'^<�0;LmS9r����7�H�͋V��΂�&%���hUr�}��ք��Q�=FmdW2Aۊg�ţ�	�`����	4dO�ه~F%�e>�i�%��Ng�p��o�V����[bX,�4y`sx�c�������ڠ����x��-	��7��T���$���$��<�`"Cn��������M��^_b=��E�ݘ�&4<z{
���Z?{�O���6x����$�ͨ<�,G���N�gp�4L��ֿ��٧��N�f�GZ����K �FP���;�׋��O_��N��)�1֦��Nm��-&�F��}_r�����W�m^P��$�~$O�(�4K��$���Z�`��y�[��֐k��J.���#�z��ͱ:�onOI {��UB$^�%s9�A͂Ү{���8��=�s�ǐp����hⵣ�jHp*�p����$�1��	M7��1Sz�b�\��&�'l��AOi٬B���B�]-��a���R��>�K������/�#�h��I/�/Xh嘤l���ِij�jhQ��ɉ��� /�Jw4�Uݭ�f!ǜN;*�s��ԁj����b��
i,u�ʃ���)�͒�-3�L����1�	�����{���ڀ�	xlgI0C����B,p��W.�c�Xb�^F��2��9�g���VG|��H�T���-��)T�x�f_R�\�R=����=��;uܬi�3���;�P��4�R�a+�nt�m���{��<c_�yF�w$���c�@mo���2�ѧ�����]P�FƕO{H���b��}��m�pS��c�XghGS��ګ���恕�rHwC��>ϻ�dK�xb�,���PY)���kh���<�R���A�cM�㵒��.���g���&O���͆��,عl�m����������2�y(`�%{�^~%�ep⵱�o��5:���d��rT>�]>�X���s��S�I�Ұ<+݋)�G63;�\|�rC�v �M�[57�)�8BH���g�����։0�J���͠�b�M�C;O�v��4�-"bf��3���#|b�㈘�����1�'���`��9-�ja�Ѿ{�	���[���^����8��g�Bw\o��@At������������ؠe����=��Trs��<����N��>�W���{���DC�皒��$ص�nsܘH�h:�ԩ�x�Ԩ�q�kvr�(�$��sqC���Mv�}H���"���P/)ݪ˦������[�g��%�rT�^5k2�L�rȻ3�P��}�r��0O�%��+S��Y
O+�����{Y_��7���6/�����CX5�LF�5VRdz��P���e���Mr�������%����t��f8t �îՀ�=��2(��tL�bc��}��Qm�ϡ"(y���-�a>,�����:4��j�
ۡfĦWp�#L\�wͥ�x���{X�_M�ӥ�6���zb�����yQ�ք�y߅�UW#1�I����[�9�Өu��Um)ZD�o5^�W��;q�.F�h�����#�� C�!>����p���\�]��k���.���\�>���{���w��N�tᦍz���=%���="ّ�	��$fH�#���[��M>�ou�>�Ҁ��_����؅�|���>Oص�q���o��-?�����+���&49����!�F��a(��,k��]����)�����Y��걑�$2�c�q�-Y�g� ¸������b4Fa˾��j��YK~p��dJ�m2e�
�KXwV>r]�X�a��c��9tv����������ͺ[�Tʥ5�!�mKSVc��պ$��۽v��8>��u�_3����j�׳k�+��N"���$C�v��4���6�G�5��B�[;*�+90}�5�������q�w���Vd��s�j8ۋW��)��oV��r����h�~r2�
:Q�q���=�1oZN�akO?Kh�CZX��F��Om7փ�X{�T�1��<[��< �ipX\c������..ؔKSK�{��7��0��es�Mh�bas�*<>��CYz}����TB�v��'�~#��4a@�ys�=�+r�h��͍�܀|R�țV�ց阔��}�M}*x5�l����G��O�8��`q�f k��j�0^l����+�8�9���0s���g�CDpT^8�#����1SK�]vm��E�P,����.�{���$�YpX��s�UKb3��"��8�Py���\G�m��Fo~�ף?��{[a_s����O��4��ʈ�'�����T�:�(0?,g��5�>frCz{����޸����X�]�a���c]�M��+��hN)Ag�e��� ��!����K�Šl�U��>����e�jV�<2����c��,��^~x}�\c�{����B�f3��x��(#T6w�0�����r<���v��*��r9���4�	ILh�i�O��v�>��<�o��m�,���v1�����[�O��&��֙����Q�y��%�e�GO��%$��*G��3�����>�Fn?+x3-�"�2�<��Goo,��1S���	P����7��1?t����M�[�ޑ:� ��61\/����5lA�'��6�N�lR�����8�O�_0,�4p�/
���i,��4��N-1&כ��a��|�]gˈ��'�=����7��}���"�ƍ�<���e����xV�g�R���
�3a��Pyq�X/Ϟ�)璲c������ ��z�;������yly �Sܜj��:�G���;���l�L|�R�A�@i�kG��y�Nw��h�-����@�36S�� ��1���M
{K������x=�>��3 �c50�ʱ6B`-n�Ѽ�����é>+�OOa|���~-���4�o�V>ƴ�PI@q=0P��gvx<��	HO����h�0�G3�!��Cx1���:"�p�n�w{�e�k���fXך`.�+�* !zx�3kz�x���C�/Y�s�̣��*�~����� 5�e�m���B��1�g���8�M�[5�0!�Q��C[���O���3��7��R���)B�O�1��Xg~�72�g��wp�@4��-�%Ԏ��	KQ���5̃�����M�-��qa٘�}���È�+�e�K]>��Lh�d��;�g*((q����r���ʢ�̭��Ӥ�r��c���$L�nLk�k����1Dyy��y*�e�_���P\< É��\F`hg{|��<Mģ��Qs�d׭���
�a�tk���[���@�SC����%P��ҥ��/&}Am��&��8=d�5���4�ZAX�����c���@��QX��/27#CdDv�+	j����ڳ^~�va��P����ڂ(ۏ��}ą�k�s�D�SLrO�>�X`�G�be_�#�<���u�fyz�����y%>��ȗ2�#�I�E)H%O�k7������=o�ë�C�/��j��HG<� ��}�<��#*���~I��̤��t�}�.�<���$�`
��%�!�բv�4���9��6,e�Lu������M�[u� ���~k#Ҷ��%R
�d���0��9!�2��{--�4)4^�������#C$�(3YhT�FhD���#I�J>�B���L[�[����K��s���	e%%��0��pD/D��ʵ pl�=������{����w�+<��3���x��_����7�!ܻwoaۗ2���},|�C
�������A�~!+�XɉV��{��/��/��w��z�-�0n�(1�H��IX���'��W��Փ`�紞�{����>�9�r�駟Λ7�\��W�b� G(����K>�(;$F�.��;�<'=���v���o�'�0�o�S����9ioւ<���u�|b���� ��ғ�@a���4�y�I/@a��x��%��9��A?��7�>�y����b����Si6%7���>tRΥ)�.�����7�M����>��t�H��	��$(m�M"Y;����B��X6!"�8��ןۂ�k�g�|NI�BJ(�K<�����l ��wiⵥ���E0���oozӛ¿����0�,�'BP��	%y^�SO=��o�&��-oQ4.�ݐݳ�>;	U�|���"�m�,��e1�&�Z�����	?�s?~�G~$�������^��;�>��O���ɟ�^�������{����������y�{��_����?���w�w��������ַ�����	�������QU,R�y
I��wm�}�>D�����6�y��@��\c1���gv��1� f�qb�y�Z��!��)#}�Y�o����m��� �.ڻ��& ��O��F�|�օ>&�&���+�kPApf��FO�!��E�F&`A]iCwH�&y�)� �/��)���1A��{ګ��p ��Wo�~J�鵕UZs@A%�K��KU�~�S�
?��?��W>��?��虳�Dp�@A����-�����<�1�Χ�D�K"��Q�3$o�[�*�{R_�/�^��׆����o~�U ���o|�
zQ6����'��Y��J����?��?�F���hx��G����R%�]��]��(+i�(S>v����~µ
y���`�b�KD��������Ψ`X)��ҫ���kS�~����ڗ��t�y#Qq6�3��x�4x~�.�<S�r	�[]c��dϟ��f�I��
�8��o0}A�~�๣'z��jfsP�~�C\l_�fv}��r=��BQ��2 ��wkh�1szu��������^;k�����b`������G>򑏄����W�*����¯��*�l�f"�K���뿮��g�gUh�p!��8|������9�b��$/��_�K��c7�<��W�R���T�g���w������u�nIV��:��������H�a`���Jx��G�W�
H�(I�"�A0�� �"` ��(���d�����S�ջv�Uo��v��3}y����>�T����k��aA�'=�I����B9 ��>��ƹ�ƺ�U�by��Nw2b� mB���n�k�&R�Ë�5�D��+���nH��5�Y|%��?:t~Dܴ�龇We�:�6��3�֛NBZ��f��m��O9������]�6����r��gOD��s��9�ί�Gd���<�J/2,lf3wV���,UwQsݹX�;wW2��Q]ܽ[��҇�ȵ�^8���� ��M �����E���%b-�(_�+@@}���,�������Q���o~�t�+]����կ��`�17p�jFu�(��e�X�>��#�p�J��9��o|#��o�f���s��X�8T;/{���կ~����>�7t� B(��v�i���PoH7�э,�W���F���GZ�/}�K�?�{n<���1��V���j?�Yr^�MLA�A���0��y��F���̆��J�#fl��%� ��ï����%N�M4V�vW-?�0���f� ��z�H�6녌-M��2;��O߄�>�T�5띺nF����9���I���d����ٌr��(�8�R�ya��B�S �M�����'|D�|���<�]$	����O �oy�[L�q��^�����g=˸�׿���V����W~�6T�iJ}(	t�� �ܠ���F\p� ��b�3p�ؤE�Q��Cu�k\��"��y�QG|g @��Փ( 6�A��a�%4?�"���?�I�"#�����Fc#O��^O��L�@�|~�F�H	`D�����4������=�tR���͕P�u��/+���,��gb���}I�wm#ws���+Φ^�%;�M�.���l�mԴ�,����żI�.���b���������M	��r|y��|(JJ�S�������rq�xXt XX���/6u�npӏP���w�����Oz��=��/[Z�������5�yMz��~����`�O}�m�B�C0�T ����w��6[��
�F=AH�	i�s�����ːB�Ҽh�a8{13Z��7�8|����\H�/�v��j~2�Z���h��/R��@֌�t��{�܇����p�ɼK�h�)+��=CX�Ս#���?���ľ_���]�W}�������c�/��U�E��!��}s�S�K٫����	��~ G0�u�����ON�y5�:9N&r,�5.�Y��,�)V5SeF����jS�>^	�7幩ܒh�ˡy�駟�������(L" � AX�<�!�Ol�R���T=묳�u{ Wp�,�\0�{x0��l�T������w��IP�@����~6��E/2��=������F�C^h#����^�����<'=�я6B��D���q�TD	tj�;E�I��	��FQ�G�CS��92�,�r�1��E�ϑ1%>/:��)�MX9���.��i�ԋ�Q�����,J��9"���	�B�:��^jt�����n[���)m�NK���iwu7M����v�t��B��o��2`o����KU�.��3U��E�~5�B���p�<|��&�2�nW�LvS硱>%ͻ��m��f�J�ő�[��%Kہ_6���IE�!������b:�Q�S.<��J�^%b��A�W����\�n:�GP�ť����K�Y�M�oL{��Q��?���J���w�{����2��j k�׎�b6O�]�*餃�L���@`{���T0P�@���
�  �q��Z���E����g���|�3V7���<��
P���Q߯���R�q��t~�����S+�����0�Xl�}����s�O��ӝ�.F��7���4WE}i]qܶ���π��t��@|��<O�a�t`�{0j�	��J�Iq\gDB��x��g:O"���������9/�DgWT��x}��9�bg�L�g[uZ� -��iw~ ո���Յ-��N����g���ݭ�d�9;%mo��]�Y��L N���v�����睊^� �Y��Rlі}�����?x��G���Nա�m�e:yy)8�KP+To��I~�c����w�fU��T�c����Rn��~��0J�8M,�F�/��3�iu��٫��㲟#��QUA�.��D:w���'�g��w�3=�q�K/z�K�]�r���/~�����ox��K_�R��h -�`O �3�i��]�;�������?m���緽�mt����|��?�3�o@���!U �����$�׸�m��.<:OKH�������A;��G}��@���ML�T(��O��4��"5N�+�{Zfi�Di�;�kIҷM�J��9�n;���4N'r�������E��R�Z'L�[Cs�{Kou"¾�>�g�z}�2��;;S�R���8���-�t���U�o���Q���~�� 4�F���\�;W'�������jZ3���<}�����_#d���v��_d�K
>�ӕ����.�W ����%��C����-o�~��϶�S��X�p�P� _ʺխne�2,a@X.8pn�"/ -�*�Þ �]0�^U��׏~��V�{��=�;��ͫcG��[��ԅ�~']�;]{��Z)CG����?��?MOz����#x���'�0�����%`.��&�Ϣ����h������xA}�I�r�β4���[�X5;i���y=�:&�vZl�<'�K.����(����!��Tk���D���F.��P2wެǕN��-T��+957�A�/�q����u���Qi ��i2D���������7����/[�P�]�,<�ϙ78^L�W���׆��/M0�	�����y�W���г��Y�?L!�-�� ,a����n���������KU�~Ŀ���oD�'d�wǾ��R�U�h���D�f���@$�������2��s��~�3��?O/	�׏�ۈ� ��?�4�֗�Du��:ʇ���U�g]��\�꠆ZgۨoG<T-���ѝc=i�-�I�ec�q���$�ɶ]�@���,�5�@��-�a�[g�w�ο���w:��Y�_m�x�ͭ:}���g�5��t��g�?p�^���V�`�m�).#"6�;/��W1{�|�>ZL��뮠_"�����-�<�2���w�qU��>����|���}߿�f�o�#�}x�=���fxr������+��T.�V@ m�u� ���Ї�9眓�����>�TD׿����	�<�����@��O~r���y��z�#���wX� Vp�t����'?���Ї>�%(�K�'�iY�N�'*��I
�])�O�D>�d������W��}�B}�<��T
�n���m�5O�y��؝�)��Z�3Od�n�7_�� ���j����N�w�
뮿/�O.�w��^v/�J�dS�����
�����y��U'���� �,�EҘ���E�}�<��e�#�g�Ӹ^c��@?���;���9�\�nx��}�������]$ .������--�p�x���- �8H�>0�Ć/�<�A2 �����>���IY"p�0�f+��q���酓}M��@* �c���ß��>�1ۨ�D��s��UN����z�3$�֐�ּ�UM?�61~~�9�8�o�Ï�gO<t�E�T����nz�E��Yq���ĸ�:��"�=�&�l�?
�ԅk�w�yP]�%�䒆}�9��,h��<m��R�8}��f-���ܹm�v�,��ovLj �rg���I]m�Fn`BU,Z�{7)��q|z��N��|�I]*��=" Q���y�w��ǉN�BwMw���C�� Z��{p�x��T 7��ҝU#H�� M�(�zzބ=?�q�zy _X =�a��!���(�CϒtU������Y�s����g��{������/>�7E}�9�˞<�8��>�o�k�練�\:rl�? F?<#@�T��/������j3�k��H����K�Zx��)&L��G�D��;=ϐ�S��L��2���G��ఖ�շg������������N�:�|��?�K����d��-��5tDg�aT�K��/����K]m�۵߲wq��=x`-��;��ͪ]X��Բ����D�W���|?Dܛ�0B�p�H�u������r�t���&'}�C�n�/�m�"P��43ɮ�YC�<�~���y9
�"ҁ�'Q�/s�=�~�ߧ-6 >A���X�-�3\D��H��h�ox2��z�ĂR���uq9}�3����x���u|��6�� ���h��R�RWbV����%ƈ�G	 �.\,lo�j�nBO���<yQ����"ǭ�)��[/�=_ש=�����{ �`��K�Z����VˬdG����[�:�h<)�� ������1���S��!�r��붽4T�u<��}(��/��u��I�媘J�0��O�9��� �G��b��U�c=y��Ɩw8���		�?r�g W�� xl�b�j�e g� �8{�X�N��q�e>|�@��"_����rK=Àv�j��B�n(�Ln,Su������-3���o�w~�Q�tt��.��D����������UNKˣGL��<�E�S.t�9�*���t�$9ɼ�qӵ�	��^9�	z`����!Ƌ~��+���.��g�������yB�|x�j3�4�_�4��آ�����y Xv��tn8P�j�2�A�����;��ݴeη2H�gv.�׸�����ù{��w�N_/��<�u���_`��Y�'�W��Q��N�s��6���d,��Ͻ8<���������?�'���uO����ׁ�0��!��� �P�@���'>�6R�����b�������q˰��%,s��7$������E���\	UtC#��F+@���o��6�x�u!�N�����~���=���fHt$��U �������;�7Q�HR��Ƀyi\��k�E�|=K����{/a��y�f=��ݙ���,9�G't��y����_�Vw�HuV��8T�:�-a'*��cҚ��*�vWst� �8t�NO2)�w��'�ئ��6����_��� :[[�:�X+/��K�d)�d� �v��1Z Q\]����n"VSu�g*����W�? ��N���=�f�P�`#�8`�o���M�?� ��[���'[�c�j�QP���L5�]���T+!��>cA�)��.�F��#��_1��t	�8H���p��_�?�7���g����<O%���T��+��|�W>��R}a+����esn��]�=~�o/�ɷ����+p0�Zt��{I��3�3�\é�>�g�� �/;��RqG.7r"�j���1�yzN���UE�9�W
Meǚ�4��m5.��&B���󗠋�D�����2����t1jZש<T]�����i����<�܀Ӈz��CWP��~���w��������Z:p�8%0�]=�5��Y�ё��zv.hQC�`�ky�m$!�㦪��;$ ���u�/<ǎ���H�O��p��>�t��ϰMd��%g�<���8⎧Yi�����p�[��oJ� �`����~�ޟ��Sm�DG������9��Se� ��Իky�ok%a��x���<2s�FwH����:��F�ߘ�����o?��J��T�@K^�^u'n�Y���(|ov�+;�`#;3�wU��o�ta9��4���_W�z#�U�XZ �P┢�kM/p�>-'�&1{p����������'&D}�'��G��#-@_��׿���}W�r�i'�W������*&����XT������>;���5�yM;��K̹��?)7u�$ҷqA8��XO�nÚlQ�����h�������YW�I���v�P�,����ӡ�Y������F�������яU������;S�[�.A_v�&}�wj>����{#BIT�in��,� �ZȆ��a�9��c���B�U=Y��y�5�g�T���%� �r�+�N_� ��_F�ԫ���YjןTL�p{�hE1�
�l{k���Z���Ɠ���F�x����ܧ�8M� ^�l�Y0D��rX�6h_����Gm��K�a��\=9u�V�eC�O�ɹ�
�����6�����.ʃ
��.��G@�ܰ��B�R�>��ǃ\�l��Mh��������	\<oւq�'񶷽-��3��~��N�����u@�hT������T �{,�<�q[��u���/}ݢy���&7$���>Z[%�d����X_?$$�o�w����u1ʻT���8�����&�������g"��1K�b�vbpA0;U���+���~��sk�랈�zӛHΚ����������C/��u�.q�I�N��O戫��e?��~��'>�R^~�G������$�V|�J\���q����|�r����e�<K��D�X�o~�`�<�@~���o.p���Ç;�s�W͔N���p�P6�a�	��k@���/��D�*��if��ZN��_���-�^�>�_�Jg���������j�_ӈ@��7�i�͹��z�����h^De�8F�&����>�����oOi�G�z����h��g�u��[-!7;ēy���=<������f����û�_�1!U���!�{	���Ҋ�_�Ef&~���%2���������D�K!�t:1�����o/G��ht�Zw+;U_MWZ8Q:��-m� !�օE@�{:q�?Lzs�v.�[ǭX��Y��\�s2�3>� }.��Z����>a��~0���w�~R��R��wu� ��@�<��ف7��v]"|��=�����7�]��zի,>�ò���'��{��}�[�j���'���nH:�
�J�^;Ks?��s�$a��]�1_?WJ��T==#�Ϣ31��.���I�J�������@7��k� ²n%��5�I汮�5�'9���[��_*�w���v? <D��#-�~^jZ|ު.�T�O˝U�>�R�?Q��8�b�C�YV����V+�ٵͳ���sǼg���t�9f�Hysh���OM����H���4[|;��~���"k�lC-��	�D���j{��>7��O4��gT:��QJ��\�,B�k|o�h�@�X')��`����J��|�ә?t�t��iV-�w��P���*�_���<6x?�o2K��}���6� �@�.������^�b7i`FT��+�V0��������J���n���i���M�8����{�2]�L�i��˧c���}?p��^6����}j�`9O_��#X�jx6bDlgÕ��b���J���﫪�'���՚��tc�y��	�ϟ��g$�r���ܢ;j�{�3:��ks�eus�K$L���7���d�\��aJ�y���m�z�䴳u��s�����Ns��W�7�|!�� ����laN�mx	�j���\�/[|ZB�0.��iU�������z��tc�Ͼ@+ˠz�`:vQ�eb+�������N�����qR�
�`�-���0wn{W�Z��ywH��2LDn�Y	hE U�N8��+���ר�i]����w��'SJ�9��}�W�El���J;����?�2,pp9��o{S���0.&�7M���=���6>������|�qj�f @�;�i��6�xF��R����$t����P��?��9� ���Df��W� bw��ݬ~�>`���Pw9��|��`J����>5&^բ�������*mF��8\_�h�G�J�2�+A�^�l>�`1n���Y��X�F)W�%3#�Ӽ��@޷�� c�<.]j���~�5���{A��s"���j�𷳕v�٥A���N�'�e���.$·{�~q�����h���5���T�I�g89��:�4�q��D"�J��z��i�z� ��������(Q���N�:���� J�g����> ������c��nY�qx��'Z{�w٫;|?�8|'����C'��.<�<+eǾl����Z�\��o	؁�E�����}���������.=�Y�L����I7��-.���/��R���tpK9�4u|J�}�%Ƶqlb5������f��D�D�4����*uq�oz��cv�'�7.1�M�J��|��bn\��	­}��~U8����B�"3�d���
�JpNT�W�;Z�ܡ1��4}&uw�G�͵~өW��끙eB
HM5Z��	�Z?l2�w|]`���6i�hah<���k~%�m/!⤴S��������}�\˲:\����~���qX���\��w�bC�:~^<�>����Hc)MǄ�A�~phkO�!|G���>ZދK"�:r��:���u�{��ݦ/o� ��cj��~.FLE��'�>.��@T����'��P����kV�Z��8c�ml`�X�ei��Z����y@n>��'�w������ϻ(�_*@��:u��Z���5���.!�g̶q����̩:��ᳯ�H�dU��`g��u>�����f6`�-��j��r����߼ov\G��j]���OΈ�Di4~��ƍt�����k�e��J�cS{.I(����S��ɧdgi�B��o}�s]��.��~�k_7P4����]�{�=�Ӆ��zw��N�=�k� ��3 u�ā�����؎Y�a���.j	��d�G����.�o�j�H�Y:�C�Q�'��?�?O���e�����7κ�2�|�>�Q��[�uN�@�38�}�1}�ވ#��^�O�2�eU���Y%Y��#��Y��,{����o l����ͣ��w{���߰�de�����;�������r����$�{��zn�y.;��N�r��j�L�׹{�f%�f��}4�5�^��)0Z�%���)
���_�<�D�t|� ��]F��>��<O�Bu� �M���;g#����2��f�T�L޽��\��f�.�P �6l�U6p��O�$]x���f7���Yۊ�a���6�Yo������~j���D�տg�I�h��^��>���g�辧u+"8=T���bf�C��ٟ8��e�clgr�nq�
N��t�٠ sٙ�o?f��/[�kz��_�3#�`���WF[�.�D�1��ͻK����\����� ��J�4�Y�s%{�`��LI
��go�y�I��� q2Q}�sO ��h������ٷK��4��lX"��O��OЧ��2�'�S=���0Y�Z�0_OtL�(��Ҿ��xJv�z���F��fi��H>�`��R.���=���3opF���<�,�V����p���yw8co��W?�����.�>N���| I]�=�S�o�'%ɠ?��H�z�q�aZ���7mD+��R�U��]�H�b�!�}>�q�����=�3�z`�8/%�U�ʗ�:θ���L|ag���Fyf��y�̾��A��o�}KT��~�E"��֙�Z �q����y����Ǡ�A��e��P���h�lJC�%E� �E��>�5 7�w N�REYT�@�Bgf�����#-��;UԹk���y)K�ćRӒ�aa��k	o�B{x�#u��`N����/Z�0� ��w����8^R�sI�0R�+��Ƹ$eD���1J�Z��i���oT���p�o� J}��,�m͇2=Gi4�������%9��f>ѭx'"��ᬪ.#0K����6��|dN���]%�Ifo�	c����R�Fm6g��l�e��d}���m�C�ӹ����α#��⓻:1=Ǥ� 	$�~�M2���:��<���{p�D��TP�D���}������J���t_�I_��S ) ��毪�� a�W��p�g�yJ��1H�KRHH�6B<:a#W�s f��m�e �Ё��_��W���.8��t�Ӯj�8og7]�%(��9�T+��_�r:�;��
��t���u�ft�Lǅ�R�tX{ck����MUW2o2�+JDx�@���5]:���r��!>�uc]���Ҭ�_S*Mp��y�uڱ�����8�*\�Ճ�\�Ne���(͖;]mkÄ��w��v�K�q���/Ϳ�V[�e��+� }X��C�i��.�=����j�S�ä�I�m���θ	=��C58B�PS	bKH)/t�-*�(��\�.7��Eu�t>}q"�F������/�}�� A.&JWj��U�Ǡ��0��`�[�H��h	���) >��#�*��(q㽶��m�6M��'P ���/x�ҵ�u-��'!�E���7���Y�;�񎦣�>�Jq:���������[��V�]�z������gӷ���t��a#j�K ���y�-��}!���M�lM'_�S�fI�����Sp�̰}щee6zN[�F�u����N�gӝ�����w�}]�Hg�M#�F�����q��v����cU�	z�������}�ȭ�*;y���Z�_��O;~tJ�LL�q��b���☶�[��A��f�n��{v�Z7�+�G�T9f}�Pױ�(C$z�2Jys�O-*��/��-�請̷!�K�٫{<�D ���3&/��]���Op�P�PB=>u��P���3��# -��Ӄ'�{�g��ǍӧT���Ї����nw�����v�|�׺fz�_��������6��������(���0��������N���7K��?7� W�?Ļ~ � `v7�E��;�7��z	T竟{U�
�j�Xr_���~�jQ	v� i=X�q=2�4�A����$�������Zpǹ l��VV��+��]��l�g.�cL������-~��G�U���� �"?Q��=�7��i6�O�$�!we%�7�膎�nP�=u�����I��[���f��	���?�rah*Z�K�#�/-�R}�(�cݮx�+���뿶���{���g�a�� @{ :8p 5�)ox�d���(\3���xG��ծf ������&@G��� `��@NJ�e �����U-�c�;��������w���� �8C Gl��q:W?���w��������@ThB�6���o��7�-e?Gt�Oq�0G�x}ε��e�<��U|�������-��~x��;����m����NM��J�[�ƕ�v)�q��KTR0vMM��&[ v����~B-]�sq�>�w*k�wAv~�7Ef٭�[5˶5�;q�m�؏���.V�qf�)\�X��Tp��#�����	v�~�1(H�Z&�������SQ3Z@�γ��K���io™���(NıE�����n�睛N9�}�/���[餃z�ӏ�Z�b�}���7��O�8���N������[�n� ��'?�~���w6 ����蹬eo6��p��pU#���U�z�t�k_�8s�~��=��{Go��G����@ �s���ԧ>�>����_��W��i����ӏ$��z����D/!L�xi~F{%n���:h=���^���gS�pX���A=�ߝՙ�)��m��Y�Ak�m�7��$:�:�����ܻ��\�ުkC��i�Us6\�؇�\����!����O�w�; ��I��aVM�i�e���W%Vy#�iDm��Fl�T��z]���;(G���#��@Y��Je�>S�����j2�,I1��}�q���B���!5�'�l�q��Ç��?�yL�*�t��S:@��~����rի�"0 �BJ ���>иup� k��ny�[f��_p�p�F���W�U\>�����C���H�c�#���>x�O:nC�	ϛ���V��	�n'��hq���̧������='͸~/A�ߗ��D����D>�t�$��0��0���}����ؑ|�d֙�Ь�G�������H��ٌ��kc6�A1]u����z'{��;�mhG-�Not���*�vC/����(_~ש{R�a�'H�yp��n7��lm����F��FT���dʨA�-�?}Y�"�>�#@����'���� m*�$��M
5��-Sk������"������0��%C���/�q�g�y��l�x�;8b@��?�@�9@��c�X�/ $p��{j�w�[���>l��"����B�+7�͛�������@����']�rWH���_���R	Ʌ1���8=��H?p�j�WP������D���礵Ou��ɪ��Ҽ�s$�Q}�="�\.�=2lP&E�,�t�z�*��z߸zU���%�|OHU�ش��b�ū���k�a��V��@�O�S�������)&� v�8��#�&�g�����U h�z�h�.�f,JN���α��O�XJܮ��{/�k�Z�拠�\8z6`ӡ�Mܝ��"�ҷ�9�/��m1V WLr -�;�}
�����=�yO����4= l+� T�����#?8=��<�� GUγ��,����g���n��|����.���׾��`O���(����?꿳{c�x&�&�4�U�L�~.8NX�+�<��G`� ��"FE�й��@I�Pb�̔��V�؛���~nz�E�=-_��^�F��	0�����[����J�r֎%����=���?�]MnM�gsu���(t1r"��m�V���mU\�bp�k�tfu;��X���t �k�N� 
/�����|�L��ᡈd6���o �ٹh�;i1O��4�k7l�V��-NN�����e.<�.8��-8l�Ӳ�Aޞ�oC�A�$SN9O&Nn�TNC�>G�_}ҫ��f_Z�_̬����������*j§�����s=��� �����Sҷ�sn��#�'�.�1Ko� ��a#��bz�3�e�_�{��K�������wB���7�i�LSN�/��~��>iZ�EH3Q3��vn�����[��S��^�*VgXe��.����i�ס��_�\:��?��Mh=СG�պn����z��9w��ۣ�;��Vc�]���ć�E�������u��7�h�O�P��W�L�u�yJ���g^t��M�s{�̈́k��@�SSݴ�ױyh�z�����j�[�ඐv����j'-���`Rf�j�jv 5�<��Z����ˬ���i���\���`�w��E��Y�7��q�ޘ���%�ϸ��;2��ͷ�7���:ރY�������~2�N,�)���Qp�8�:�<��
�T��Q��+�sę�����4JR��r ����o��m��u�Y�==}�����=���PС���!���������'�V�jDy����;� �l�C`�W@:���p�;��%ԑ^6��<��R	������c�\R�Ui-�����SR'�k������VH0J"��~|����g�G�8~4'>��
�h�Y�:=�`N��V~S~��s��.)NFa_gA"��d�D�pG��9UXK_��ˬ�}�Žt&9]p�0ȍ���Me�⪘�gS�k�4_�{*D�4o_V	`J��0���� 妪y��l���[%F�eO`�q�
hD��\���;\xq�
?�L�P~�_lw��Ad�W���Q/�5$ZA"�Z�x�s�k��O��q`����<ň�?�q���`)��TB�������T���&:~�c��ϧ��>Ϩi�~�FeL�_2]Zw��<��[���m��g��[vi m��Jх����|��y�r6��J�?$���kKC_51_�@?��L#q��k�ʛ6S��8��ꓙ��0�9��xZ~4�x7����.T�R[�����n��	��'X_�E\�^j��6��|�	��F-8p �9+k9c�?���K�l�7�)����0-�cH��EN�~�����E-��`��Np���Q����&�J<1�ۿx��Dϑ�>xw�k^�$������.��·㑮�@G�����g4��V�,i<�u�r�?ơz2��I�<f����tslA����l����)#r�"����T��	���A�m�m��o�$���驚��O���~�s�0_d���{Z�����Mv|N�w��\�q������l2��sY����^�M����7��+(i��p�iJq��� K�(/.��;�1P�����������3r�T��r{	 \b!\q�CX8m	 �b��%Ps� *&�r�jG�r�Y����/��/��&7�Iz�ӟ޻�F�~�����T���^��h�\e~^���+ш��3�c��_%��Qz��{5X@�����  ՖI ����ц�Z�$�I��V�����X�7n!0g�?��0����� /d��U�Qp"þ���P�������]́�
�W��i�E"�߳;�ƕB�k������K
��)���+��"�z����^�.�����(�DD�ʧ�n�c�K�G����4� ��s�����x��C�.*�1@̓�����luA-'w���$�r��I*��U���>wp0��@�؉��r�u���q�`��/?F�=�iR�Qy�;��S�4}پ~:��='_o����X���Ҥ��Πv��mf<m-�}%�APbUb��@�&��D�}uÐ�N�I	��il�$���|	X&�}�r�?K�;�5ݕ��)+�Y,�.n엜�u�)��E��=6q�4�R�K�T�)n�D�T6S\�J6��g� �`	���4��3��:Ϩ&��)T��B��u�}��p!:M��L�4m 1��б�7��I\�[���!�V��د@|���6aO ���  ?��6m���m���� �����8�q��J�_$U�6xK\��U�z+����T�������2��j����&9�d6�S��f���o�;tq?n�צ�7�
+��^��n���D	�$3��E�l𻓪N��-�K�7���,��K��`Y�<��p-�< �].�I]^�YZ/)7.`-<U��Yg5�d���z�F��@����dg���8��h�Y����Rv 4���`�K�o��#��Zvqx盞�s���u���!/f�ʈ����&+����i���ŸK�|�B:<�Z
:{���;H	H)�����4�@��m����TW%���'�"P�q#F�ƞ�>9�^2VK�h�h|���l�u���O�QSXb�^�����W�v.5��te�;u�}�!���D���U&Ŷ&��.i�G�~>���q��H�V�(���sr�\�� M.N�����R�6������c��\&}�oL[�ο���c�=�����Κ����@� AΎq��Q%=1�������DD�/.o��iU���2��aM�o��O�"p�� ��p���Jw�r���1Ɣ��A�O�~�)n����V	�:�pp���	x�t8u˃`<IK�Ƣ��L}�� Н���}�k#���)J?����˲���t�0S:�5z0�;��P���w�U f��9�< �Jvl����ܼ���|ּusn3���f-�D˔�hU�oW[�c�G;���yй��W�ދ�Vuw2�g�Z�6�q�����df��DPw;���CV���Kd�4|Wt�%P0P���#jp����
��'���5�n�h��V~j<��A� �uѺ:%��ߨL��%�k�~�����ۋ!����<���KD���v���S 26L��A����kD�w�k����(T���&�7�Lf���o��#O����4���s��wZ� P�䁉���ȕ�T�~�!��t�l	��������d\�k;��^�=l�����2��R$�h��s�w�L����ֻ2�-$�F�h�M�|˝�m�!�D� -�:�J l6��a#̪����"�qh����%�
�yN���>�+���:� �j'�#�����Yf��y�бɶe���N��-S�q|��E�1�r�%qU�O��	�q�<�s��6��A|z��	�T�S��ˣ�#���'N�{n�����9U:x�������;6d�R����^3�����F*\9c��/|�����3?�3fc�{�;��/����P�s�9v�K�2�t���o��~>/�/�q��F��o
���|�j��5-�k;<��<�t�=#%���U�g9}�hM�������϶:H2��׷�����KGX6&���^���u�5er�a_7r9����h�4�9��dq��f��G�m
&{n��J�<��Z�(�|=�{��X��S\wD���B�Ĭ����O 38�O|����s�H�.�Mq���%)���� կ����@PѰZ�@
@�Ç�c��~�Z��n`j ����x �p�!$���u��m�$��������]�+0�*q�ѺдS�����m"PQz����D���DJ׳�g�	g�}�*�=L3 �vG��,w�,:3q5W�C��q�f��k�/����V�c��]Ұ������z+PEZN�w[1}Y�[Ju���E�NZv�|�0��f���:Sd�x���>v�ͺ�%Z
�%N����Z��b�d��e�gSܠ���D����ˇ?�asÀN���m����}���~�z~�E�ϗ��%6�����;p� x���Z��&*�, �6?�S?e�<.:�wH8����:����o/OsM��ᾁNb���W8G�/��\@x�;'7�@U��է�Y9�҆�g^4�����%j��������{i�yc�{�K���z��)��7��>����w/��]���V���{>DW�ש�9��4^�����p�u����MY�o�wN?��98MO1�>�A'q�<>]��q�	W�H��r3�ߕ�+q^Xk��K���&��-��B�{�:x����"t��Eu�sp���qg, �~� Rp�=;8 5@�Ɂ!� $��㏦�擾�p�-�����"c�mz���l�ҩ�7l!pz{q��p4>ʝ�Zt�6V�q���~��>c��A����#�"j�7���K�g1�z��ڽ���u�ϭ�烪I�`k���5G��"yW�*��Z�{̣E"�k����V����c���:Q�8���8��w���t�H�!��ƅ�4���P�xN�`\o6��W4n��{TvT�M�:����}��O��q��!yH�� Ҹ�
q��Q�d ��!&�:n���ҕ�d�!n�<�6t�/zы,-T?u�|�i$ǃ.t��������9�Y�E�ߜ%뗈������Q���^g?��������k������(��^"���s�]:8rL��i-솽�4�C��4��o�u���*�nT5Su��w�i�o�� "X�4��gl*=��Ñ���d�
�xUs	���F-�a���Mj~�&�����YZ�������e]��ۡ���{:�z��-M�d��������ӣ��t����6_��)���`W���O?����i�� (�(��(�xH���Y	��S�-!a;�w�O >��s�W瑚�@�Pk>��%�x&!�B��r?��H��$q��K�~�M�i�I�Ý�IϞab{}������*����y�u�ؔ�8"����3,���ͪ7.0���F�)df��c�w���*��?�;����o�𤕙�/�'���WH��/���
׻�u�]n�̪�����K��p��*�JՂ�.ġEj�Nʋ�X;(ˋ����j��|'-k�c��ǡ����wNi�A7v���m��U�V���L�<'�����E;�dv�ǘO�%s�<�#���HZ$E�z������qazfaA�;oǯD�_��8�x�l�I ��Y�y��
@X��>�~q0�x�:�g�rt/�6�ܐEyx������|����A�j�#u�B�w��1f:5�T5��tӱ�q�笛|�;g:ط���r9W�ߪ�a]�6Bo�P�,�;��*2�ft����<Q�����i��Z����븽�&�i�%���#��I��������w(ͫ�t!��5�j�g��˪�t��f ���{Ussr�P�%����ެ�
 <�*��v\��8�bT}0-w�z���ĩx����aH(��N�e�}����Q1v4�*9d�q2U&&�z��F��	BN�ZW�0.D/JzN?ҳ��(Il��%p׸�xI>�'&Zg�J`�*����ׯ*���]:\#�oM3�f��� %8G�эnd�������,$�up9:��iY:��j����X |��(�=���DN�b��Qi>�|}�����-N<�n
�H������敪JyN�*%A��%�'��>�U+:M�����6ݍ8����
y̌`?`ՕS7�)�n�����f�>�\�����D����sx��&�Ģ����{�K�%&�~y����,�D���%Q��&8{�LDP�k�{lz����}}R̞������D0�K\|���4�.���Ļi���ܣ| �Y�~�K_jj����߷g��@`�KX䀻'P�><[�=<[��n�J���A����!��(M�-:��c׾�}���c�rg���w�	{q���%M�D����ϭ3��]����)q��M�o�}Z��$-oSɬLC\hҠf.c���N��u����T�G��\��o��E�9Gtp>��]�rF����:�:�JK}֭4���i����|��bn��Q��3o��	�6�gQ��Eu�@���Z��l�� z�����&>|xd,��  N�!p�H�,���#���Q6�=�/�{ ;UF<S��4�-ʨKױ�g\:�;���@��s������c<%�i(I��=Q�%�b��(I8~��}�jL�;��Z�6���t{Z�*�g5u��r5��e��F3ì�x6�>��܅��8a_��7��<p:w��1Ot�LG'EU���q��sX�;��e�;�P�e:L\���6[�Z��}�esX�GÍ/�|�Kd}�X���N�HG�4<7�s�K�PZ�!�- ����͇�b���/�9�E�p���O}� �� pl�~���m������ �M`�����9O�>$
�K���ڡ�O�������^��u�jE���x�,1�\�������i�Y�AiL�:x��A?jgD��
��z�zY��n���w�Ϋ|��|���m�3���Ţ;��tP�����b�-���8���a�vw�!�v-�,U����%	����L�'�d�m�̹����A�w��>�W�1݈S.�I
T����A�;�C7�J��-�������T��	Q���n���jS)ߩ:k|^.B��)�x������t�{��\&<�	O�+���g�X�9&�A/Ї[\���g>�|ۃ �}2�ȅy'|�����3ϴ�\x�= �d��d���7+	�ʥG�l��f.q��րB�i��u�3;�����ɉ懮��ێ�~z&���tJ,ٟ^J�u�4���Ts��c�`�3~^I^��)�f�.����;G��Rc��{��5���l�3���o�Π��[)K \0v�������iZ���r���6Bp��5'
�J���n?:֣	qJX�@uҬV렻	�5Lq�{�?Ł�E�װ��\�ey�h�<"�zu 7%.��=�8<�3� ��nw��\�����]�wh��\,�=�{X!
��җ�d��P
�/Z�{���� 9Qm����%?n<�O4oo��w�#.[环��7$����<�R���޿M5H���,`���;��{?7�F1`7����.�M)Y�Z�m��}�]��eЧ��k�oJ��9hRd~'�A8��Sۑ�[5I��T/tj����܂�F�!��~9�O����_������>��)D�v*���R���N�*����"������/�}�\���6�x��t��KTh�C�w���Ϳ=@>x�H���@��s�}� >�"Y���\���e��y��r�Q���F��I�^��sB���U��G�T��qж����5�b�V���W�wl�|6����NB褽U3h8�*�`"Ɗ ߝh���XT�<}��� �t\���N6�w�x �|� �Z66\88-ג߶ӗFp����P�{�x��!�Y�V����@�Uj0=,�w,��������t�F��Y�^�(���2�_��ޢ�}���h�<�q��Մ�j���J���2�=`�ik��9@ :�r�LV�'P��#w���D���(��#|���x�r0���YOH ��ز���G�ܧоV���e�q�y>�}�����3K�'���/�=����?w�y�2Jf�̏�\7"H$��6%����q^���6�m�W�Jl��N���0d�5Nw�|*�ӷێs�s]�Y���nQG}�(k�����.~���P�h*#F�"�l�`q�p��;x���YTj�Ƈn򯖝�f�b��Y���I(|Uל|�n��-
J@�q�;/zg(qå8��*qV�����򼘫\��S� �ߞ�S���ד��a��1N=<��� �TӐ  �-���*��G^4}=x��}�XZ�����#�ry	�LϠxi{HC04�)*�i����zCA��i��s�^��@��h���O_�C���VZw��̷ݏ�'v���LRPG{'k���j�����^ʫ�|��t�R�5U�F�h�.n�W�������%wb�G�5���5o������bU\���<���l7y햭U�Y�Bں����.�z�%�1� k��MN|��z"p<��EeDu��iz�����K$��3xP�n�.`B��8��M�7����������=Z}�C2 ��*�/��l�	� SJhé��vk<�ȽJ0������6����AB:�E�A=�(�D ���0�cԧ����LJ�}�A�Wt���b4�}�=A��_���{O "�1EH�>�N�lf7��e|�V~��79�ihV=s	���)�lu�����{:Z�_���L���V��Z���K������G��h"d� Ψ�@�|�X+�m��o�YJ�x�wv��$d=R�*��]���M�����Ji/��Л ���zk���w<Q����64ΰ�0~�_4����ln�ۛy��뿚i&@�>�����~w�ɟ�I�!�:Eޒ�VQ�Ɂ#��	��7��Ԓ�H�:���oM�zի��3�;�����'=)}��O����$������׸�1�.YGy)�u/�P��ұT�6O���S"�I���S��"�P�8S��u�y��^�����z9���le8l�:��ղ���w��˛꓁w��M���\�Ra��;M�nv�ԓ��&
�q��\5פ�����lim����|;��k��6��-���%�t�E�; �xth{�灯���5DD4"^���"�DR��[��w�R,U���Uˁ��`E�?�[�e�8up��_�|�k>��ӍP ���H����|i�C�	}�쥯�@�$��H�Z�pcz���� �)�N7�8;�S÷��m��o~s˗~~���v4�6�)j����x���oz���9�(-��,��ey�����Q�:�{��9��&�����a�:K�Ձ������b����`�'L��~O�I'(��u��Ieaw�4��hDeW�J�V�5�I���V�Y35]���q-��3��m�yGqJ�HI��g����������Չϸ���w�î,���և�\/L�� ��jQ' )\,���=�'�{��v�]��T)�S$p���\yB��3��?���Q_���oxC3�����yD	D����&`�yx��%|)��_C���8��H4�\�1<�GD�]��������^$��oG���6��Cxwݛ�֋�UV?�fc�ݾ_�t��W3���x����}�av�qQ�"(`[p�0_��QnЪ;����1����ew;V�߳�IqA}�Nԋ:���\�q��vn⒢8�寗�b�E�6�Ug���{�d]%p���f7�Y�Cv����
n~�y������[�{���g?W��к��{m?���7H�_x��g��!/cq¥.���O}�=�D���=�y�F��f̞s�ֈ�KSs���t�ժū�6__m�Ɖ�z�=��F�D�$q��L���m �X�������s���ڞ�;�2tn������D���k��D�}�DE��Ş��n���MA���$x�t�9�h���[��8���&sT����M�?�x������%њyG��r���� �L�������j�M���hyC@�-��ؑ/�e�ݹ���m���(�P _�x� ]��ُ4��D�|a������ϙ~�yx��'!�-
���*m��+��K�A��"f%�]۬���ڶO�).[CI�����u1X���cSk#s���e�5��O�G�;Z���u5��}��L��=���|<����o��]Ͷ_��4_�:J����L�e�����i8��mg\��"-w�%�M>�m���<իva�;���e��z�S��-g�P�V�7����be@3\>����Y��M�2��x<���9�9)�g[�9U��jN���'�����a�1SM!��/,օ����E�q|:�|�s�����3�o�!p�pŸ+;�遲3�ChZ	���_��m�b3n�U��}�+��ۋlU�9�}��u��o��v|�����~�Й�%ǏkA̸a��ê�)OyJ���y����(S�>W{so��s@����4��I���Aǘ ��b]��;���,羮�����չ�H���N�G��ǖ�w�ߣ�����f�j+��k�e+�u���i+f�e;wR�i��b��<��7γϨ��s�j�cs��Щi9?����vnUu���G`��.$�v�¹~KH�͎�#m��;��g��t���]�^��n�|��ފ�{��������2F\��v�GU��������K���
��|�	E`�k6���s�H��s�/�dy�Yg�'?�ɶщz�&�p��t�?hEsG�W����ýt�2 �xPfّT�`�U����o�	��=X���.|�����W0�yp���y�:���h	���}�{�_��t��g��@I������(s��������m�/ӏ������ϑhe*��GDP� ��V�Ѷ��Ѽ�>��ÆM�n���O�V��;ۋ���i�1�ՠ��6����N?�����F���av��RMfͿ�A��m���ʈL��ԩ��Y����'@���ɥ_HL��Q��#���a�A�:�||�HZ��1�6N-L�xJy�w I ;Tp��F�7T(0ӄ��
��Z׺�}� ���������w�[ߺW�O �ڬ�ݞ���OQG/<�|���`Ɔ�Ӟ�4�$�^���7PZ&�e�����>�i��xG�F�0f�������:&:W=C�������\�����ݯe�
�$\*]k</}�>����%�2Wـ#uU��U��}��}������;�h�(�%��F.���=�Y�ҊTkڵ�8�i��R��Oc1���9<�W�Ճ�^&����C�Oc�O��Q�p*�*1�4��v/ ��G\_���|�Z��#�Hz�ӟ��t�;�?�9�1��������^�:S���_���I�i���������6�u
}��׹���>��6���x�
��¦.9tޮ���t�����;���׼���׏�a�D�G\^�q�⪕+�$�����_d�I���_�H��4�5�W])����^���t7���6k{��e�����R nY�A�}�
�GMn�:.e�t��+�s���uV]˳&i�0ߜW���5���ܘʉ�c6�iA�X�}g9��@�&�^9�Q7����(Mf]>�)"�O�ش@�>�օ X���}h���A>�<b����<����}��w0�D~�X2�ӝ�/{/�T�M�O��$�������c7��ͬN���+^р�P>.}�R,����hz�3�a�,���;~�^�y�I����=�BA�↨?�yVb
"�(b��<T��O�<#	| :]�7.f�r����f���C��5b����XX���KiO���}=��u�O���<��D��� D@��%�z�8��iY�T�4�o�����mܖ���N�o�N�"���P�ڿ��=G�ݷ�"9�����L�b��Z )t� C���l��$.�EM��y�����Ӷ���d��%�L�ɲ��!M@-�Y 8�F hӅ3��$. ��Q@^ ^ T����׽�r���u�}��XES>~�c8?��h��Z�mZk��j�Q�8�Қ�I�Q���e@=-yS�Y�/Gm�Z��[~Y�%ͦiz��!kM.��2vwz�fi7�d�9�RVi>D4F��y��|}��`�FW%��h�:_���z�����uKv�~�h(�w:�"n���zE�O��ګ�Q*ۇ�rj{I�u�u�	�Âp�~�} OzԤ�#�)�V�J���/Q��cP����t��A9��	�(R	����?��Da����|�.`��-o��s��X;p~ ����A�x�$�� �<n���P���}��ퟕ$�h�#F�$�E�A)O�Hq��)}����!���ݮ[�n.��q�J�=��ǚ7�A'�"C�tG���|�����n��*_cܖ�����D�}?��m��wo4��p��eOt��������ur���b�?9c.������I���u��U�Ї��v�$Χ/q���k���/J�����ϻnimþ!��+
i�	��Yy�!�AD�|e~��׃���B/���! !�n���[�~6xy�"-�Pwlc/ y����}���E�*"ħzi(mD��d��������*bTJ�@7~����i�����}��$��<��_}?���i{�EM�/�oU�ޱ��5c%�$`��/W
��O�������\�E��9��4���%7f��Ţ�WGgw�����c��lX �T��>vj�i6��牱�O��n��"�{n@'� �xʭ{��9�n"2�nh�_D��}� j˭�t���g�Z�(����*�izB�gt�j?������'��;ڌ�̋z~|#���g���,��mq@<l*#���iO�~��l.�=�C� �{h��O�"�OI�X�Pǒg��SM���WJ3:'��������������#� ��z��;�<Ԣ�si�G���+��� )��u�8���1�=m~m帻M�@U�\�[��qoVm=�f=����vwU�r�
�L���^-@3��{�+úU��q����VU�vfVY��OT����Z]*u�W~ݤ���k;������.~�ݑ{�؎���*h������ݾ��)�8�(�爦@qS�т�DԨN1�C��/C��R��"��%����MY*����m@`ϴ�΍QJ\�<<Ņɼ�2�,��4b�S��V$B��!���01Ezp��� ��o�EZ�	�($��u�
���%F`��°�M��|�\���D���1����\��^槯���>�LQ������u���̇�!5�E;���ͫ���w�ܮ�{z�ډ�
� r!L�ǾΗ,ޛ��m��`���V�oз<m���;�Ug���$����	�!O�������ϰ	��">bS*�t16di13M���N�q��܋�ڇ�b	�(�)��8uѓ0=mߑ�!�"w�O�3�nZ�P�b~��J�K�	���'�Ү߹��@c1�иW��80 ?\B#?�i��:��#?��=����� <]���mȋܝ��Ώhlz��4?�1��\Su�s��*��8Z��l<����9~��n�G�ˡ���ޮI���צ$b@l��X�϶�l�J�A�x�@����v��OJ'*컗M�?`��0��?S�u+�k�_<(��io撾���t��"�8ږ� ����mN�ʱ������/�)�T"D70?�!7^��~���c&k���5�80{�#i��k^��ӿ�u��8�������?����o~3=�Q�2 ~��_n�A7��M��UNOr� 
��ԧ�{����w���l�7�||��hG�����>� sNx�D=�x7a�	�}�7@5�} >�5~��Q'�<��@������l
~#� ?�4����m���S�f`�K��E���?E��zN1���v6�n��j9��$>���T-w�mk��z��I�=��~�H;a����mQ�%O%3��ݩ\X�ԃ���I�'�n�Pl@����w�A���G�!��vT5ˉ�}{7q.�Mp?	K�{�������B��Ґ��wUꇈ���7H3K�p��<����;����+�/�S�M��r��� |X��9���~����
�J
��P�^4q���aR��y�5ۉ� �����^�; �t T��{�g�����-����7�}��<�1镯|���w�a�j��@��L1,�/�S*��_Z4�|:oAS��KyF����oD��R�I
�Z���س��`Rv�*q6RMշ��=�'s�=��]�1��6;�;����%��G��(ެ�������2�n @ָ�.�ƕ��٬&�ɨ��&��M�H�h��Ӵ{f�gO�dƋʋ����^G�'@�s��\���'��� Z~�qz�� ��apF:2�@����T$����3ҁ � 7L`��k�U�r��{&����ބ���kӃH���w6N$q1���g�i�Ç[���@]��}�P����xFϧ$�)@�Ri�����E�;��$�ޕ�ה�oG���w��6�u�N�r���}����Ԉ�c?V%܈�!M�}Zd�/F�w�kC�wP��\;�;����߳؋AF	���np��s&��>^\� rFi��r�F~F�j��}���7����������H��7e0op���;�A��. �����׾��v�
�$�yBJ �"�?��?�g?���:v���P�<�!I��խ� ,:�?|ǉ��u���O~Ҭq��p�m���� ��mo�z���w�KT�*7y(po/>�OɅ�z�x�_���g��f��Po�)ɔƋ��}�x��?o���P�"H=� ����u�:y�.12�����^ϸ�=#^G�F�U�i��Ҫ�5�D_�4�ERw�V5�4�wX�s��"�ûM��}s� �<qcγ�p�[��h����4��U�1�F�f��������M�OV~/�Z�	�^���s�ĸޜ���vxNC�{
Q=6�)����9N�>���Mg�q��d�s�_���F �ড�G 8C����O��$�//,W�T*��t&v i��j7[f�^�y�x��q�okAu��;��ʣ��� �0�s�u@;�2z��hn@����>�A������у�g>�[g�ҹ�(D��[��^���B�I���SA���i�_��{����Ǌ����7i��ۙq���k��΃t.��`
L����y!׏�{�k7v�N_�..��}�e��uN�[?C'4��r��>��ř�}�4���z�|��]\���s�	���<���V���G7�ͼ��S�[��ɪ]��������V+m�g�81lCSu�P;�����1q�~�W#�F��	3"ti�ؑ�T�F�V��Vn�?Wi����A�M �\M$Y���u��9 �p70�ZD�EI RO�H�~9��X�P�@�C�y ��7L<C}@DnzӛZ����OX^���� u�e/���'?�p�@�G����\�n �C�w��Q6-r@Ƞ��➁��$)zF�f�x�6�lo��f�N�Pc�����^�:�t���44�&�ߢsK�+`��y��y�/"�g\�Q�ddY˜v-/f��s�{�����T�|�t����Ķ�S3D��ց4o���[i�ˮMͅi�j��٩��u:t�v����c�m�ܲ������BR���KXr��������ڹ~R��Ӊ
�j�����	����O�j ګ6-��ߪ��TK����܀u�M��;!���Ñ���8�f�y�o�q}���qؾ��6a�4Sq#О��#i������g�3�������t一&�H]����+������sj�.�<�яN��׽�9�� ��������,S�hPw�\<�z�e�mp�P� @Ǜ��&q�P|G�o��`���u������'��;��TA�����3��	b�(�>�}q��<"�@���Jy{	*�r���;S �5��J���Kӓ�[	CW庭2+�V]5�ە]�4�;��s�1���_�1���K��)���c�������h����渹j)�sgԤ5���K���o�X|ʝ<��,?��?��ɠ�������>��^E���F���}J��[IL�m/D��- �X�@N�X< K 66w���x( X�'n��r� p����\:�y�-P���3��h����G9t��:����!�X�`xF�At͌t�B��t����6��t�?�ɓ���}�z˯h,t�y�w)L�ݽ���'e�_���V������)�����$}��)�E^�,i�����ԍ}_lAҁ{�اA-����wmq��i�K�S\K��G��W
(�Z�ܠ����T����tn���:�����^��l��&����Q)uipJ�Z�
Jܰ�M܏�+-ֽpm�$�_�Fq���S�\�i��@S�P?���*���-S� `��� �D�N�� �� Sp� p��<����F|��5�qzM�����wS!���C��,���y�
�G�p�Mc����v~����|_�8}������)ŉ���S�D�n)-�
Hgi�h����Q��2��tj�C^�{�zY�e�i�]�����^�P��jP�:������q3������}<T>[��j���z
�G=p���	�b�%*"��jk�g�^C�d^gʹ�L�b=z_�HL��}���$*c�3�kZ
���Ƨ�Қ�K��� V�=0�+��ϡ��{��Sp���j\3�/�� �� �����t��A<n��,�}�[�b��n����`]�P��`��=�7���@�(�]�z�����}ﳃc�:p��o��o�Z��H�k��kv�/�.����@@���>�Ȼ ������ё��M��o����L�lb��ּ�"�h2-a偤�^QTV�410��Bg�^��>�p����u(5;��*~��B����/���]n���c�F{���>��]��ϟh &5O>Z�yS5�\r�����u��C��#��#?��M7*Z��j>��gtay�0K��{Y5^i�GB��q#�$���-0߆uQu�m:���ǆ����HCG@ �%�//}�K-.��T��l���w���-[���t��Y�w�kc;Pӂ
UJ s
^�w������"�t� �MJp��K��8�]F`*&����`��h3��	���>����}���*郣1�$��xG����M����k��a��#�yP30joZo���Ԧ�X6���<�D.^|]�q�G�z�(�>%)]ܰ���O����x`�@o�f����~��k�AfFo��|H"w�K;��Zu�1;�P�6��*��ɐ��x�����y����t͏�<X�P7#�����RY��/��Q�M�O��|��~�����n�gn�������� �Q7�X�m�?�A�yr b𲗽̸nx�Իj�Mc��t܄���7�q��>`�pr��L�n|Ax�6�|��Pw�	���-�wCR�<�����~�9���x��^:�O4���(������>�:��n"�=QY��nk{Ӄpn?�z�}�TS�:�;�s�X,VˎXe]�-l�V���[�����0�b��p_����=��������ŵln�#��q����x���ኪ �lvkJ3�ӌ@���l1��X��im��ߓH�	3��ǦpS9��G������/-�l�c��B	��{��[� ���y��@��[��Ƣ#6��E�����'uia�? 7$p�t�n`�t��ۯ�� �N��,{p��P.=o�e.�����q@@8I� ]����܋�s�M/B'q�.@Q	N��_o���fI���T�(�ߦ���1Ds���b^P��5�I�-���|?��4&`�˟u&ϫЫ�U{�.x���_u^5p�;�]����n�Je�t|����:}t�,_��`��m�.�&��ܰu�n����gf��r, �����L�9횿k����|�F���C�{]<{�49����7�	���iƛ��x��dJlA���p>?�A]	��[=�����S�裼9Ax���������>tÌeDܗ^J��Ҧ��Kk���?�����?��	�=�.ؼE �S�G����������r��* ,t� k^G�C_j��O8e�U���6�H��	���~A> nr���9�K�F�
3^�N5-���Ӌ�9�h��c�6�j�T�#I�K��s����c��~�f�<7@;{�ja�����b�Gk��w��O��鍗f��t������.��S���sl�6y��bw�@�;�;2��I��ۚ���?�{Gz�����$�;��0t�l4�G�/Hco�6p�c�vuYg�c�����Iu`;�e:6Z(&6c!`���@�k=o�z̴m��$����MP͓�J4�g�o����է���O�=2�櫜�9v������R��;�p��i	���<9G 8�c���,	��'��9�<fb�^2	ftь� Ⱦ�x9;]#� ���F2�o
���tR
oS.X�S��s�ј��a|ϑF�_;~.(��A��~�*ш桶M7u�Z/�3�:��Hr��r���l�v�}:J ��iW��ݡ2#t�\S�M������� �p@�LV�Ȱ�^6���WBy���O�,T�T����Š�h�_�`.�X3�Or��Ā`�+puX8����u[��i��~(%�YG�=�N�U�X�g%.ڿ��Խ	�,[U6�3��{�{ڃ�v��v��!�ӏЂ�Q�C�CT�PB�PdP$P� AEBCp � 0�V'��t+�/��{�9U�����e~�j��SD�}�DU����a��O1�"�P�{Џ#�b�
#���럋�Q����f�[r��;��J����'% (���P&�a�7ʠ)&��@�Y�:P:��sT�;]��j��3J��=&uM@)L]%���u�<���x���;�ى�D�u~�11�w�u=���y���Zun�"Z�~ev���W瞯�����Pd����Vn��,���b�����"i���*3��s�q���?��q��9v7�
�q�3��s��G�|"w��`�C�S�vc@N���y[������i�:��r}$1o�Ss��Ց��;�:QK@]�ѭ��鴬ݛl�Nun����G��O�4'��}������N P��i��}�i���ȇ=��=7ˡ
��Mb�*��o��oM�?��w���'6wqD�9�	���資�p�|\cE�O��3�
	�VH�N�<�s��>�~��+�8:���<�򼊯�����yC���s�n�f��	� w��mC�m��	�i	h�_f3l�gu ��ts�>2�.x�]�����4c�}���3��{����_"�u[��@��V˚������	�|tvbA���^�*�])�[;)}f��k��>ѧM�w��iޓ�[�c����N��~a��7�1�J#U��<t��8?^�ɤ��OO <1-=���T��}���8�\PNgi
 SF�³t��q�/L��O���kx愳3<����>���w~�wl3Ͻ�-oI/}�KMϏ=��Q��J����7�!=����Q�`G�oX�}�=�v��H >p1B��e����5�2�>��8�(Es.�u\#�����;�|g�H���)S�SG��L�W��:�ZDh<Q��7���>|��	=�XY���M_�zYٿ�d�uq�4]=�5�;F����>6��zs=�TGw��1n��7cl�cn�� ���Hj=H&ތ�|o2.2aj������M5��0�i�ͤuo�M�E=��l�.R��zG�0�O~>V�D�X��%�[��{N��y-g.o >�8H-[��W�^͋�r�%N��&@.���s�!��7��*��p��<�Y'�� �qJf���a%�=T=<�2 u� o:R�F,����CJy���n暴$R D��S�� 2������*��;�����տ?]1+!W��j�gQ*��C�f=������y��"�f�L�O��D�x���:˿^�"\�k�,�U��J��U���d����5�~����,�{H����?^��uTh�rpH��&�_I'���n��l[�ݲ?#Ww�5�mz�Y�9��=8�[ľ<�@�w�J�m����"PA��>�W������$'8mk,*<qQ��>)��>��/�*;��FN6�8���'?9=��5�x�����e���x����<�6^�V>��T��`@f�5LB�e���<�!��,p�\, �����y 7N
���k'���G��4�� J�/_N�zԣ� Vp�sN�A+!���w�P�qS]xD ���ϧh��$�~FR����_��� ^�S��1E�
�괕�H��ۘ��+�Gӷ��]*��?p�i��;�Cqxgc���ϦR25�or�ù�����81�o�����˷���HDu�X����UX|g����)p�r�����8���l`�`q2rL��҂���Ӊ _���b>*:}*��Y��Z�D�RD}ޞ{�@_UJ^OI�X�����V�@��r:;���8���.@�R�� R�j@0��S`�iN@����K��=N��:�p�ς� ��A �w����X��@7Ϻ�ʯ���m���jA^Ou�9�nV�Gz%�R��n�{��u͓sF�����"�g?��w�������I��(F��o��+���g�<�:�Һ7�<�L�H>$葪?ĕ���A�G$�W:�F�҅�w�z��O��[r���E������o�`�c�D���3�؝��z��>��0���f9t�r�v�},����n��MD���������X]H��Y���?�[/�=ݼ�CZ�6�g8M�iz��<��e��d��]�m]~v�����K�A�"�Nv�+��V/:i�h(d˒�O ھ/6�}����FW��b{ԟ�h1�O.gJhקY\�z��Я��Y��/�a\����_<Q�{o�g�d���>h�7��n�pi@[w|�"zr��A^���9v�-��@q�������(y�/8y�V��?}��Aesc���m� ���}����}F��`���y�M0:'��>���]	�槠�%A�����u�2,&%��͍�����A�Y_���Z�[�����3����ǰ��]���3Xt��Jh��C�k���˼�9Y��G�+]\�+]��O��^�0���v���_U��q�ʇ��ḓ&?tkZ^=K��9Z���]W�2���tP�~̩88����I25��ۂ��մ�?{m���|�^�����֠<���
�ڡn"VG\rD��E\�8tG�xn��[�"�ڤ�)pD\J���h���p� u�}�s�ucS>j � ~X�@���W�ڀ�8>�S/}��Ǳ1����6WA0�0�2}���ՃO����MSMn��7$����/�oT��\�~cu �/�x ׯ��� |?.~���dk^���/R!��=F�)3�s��o��%�]ey�U�+�G��g��r=�e��bH̓�ɴ��n>;�vc�	��T�̗��$�^������ѷn7�~��Gu����r��A6��%�� }p�<6��_����l/�`=�8��p��f�
���)�I?��<J&e|�_�����K���Y�w�M�`)'q��,��cO΍� �~�����i���Y w�9� �� �t�������tZF���� ��y(
��H����� h\�_l�#n/���Wl��[&�>���F-�w��S��z���0I��q�m�~�/��/Y9���ƱRa� =G<�t�Dsp��1W���y�|/y����\zǷk�v�{�������$'���oM�],G�΄9�$DN�;%cL�M�r���׺�������y�!9�7�F��?�xN}�=w;�1�V�J�9M�ċ8!��sM��,�_���q��{%�������D ���Ŕ���l��s�ոi���&T* P 6�� ���� �M��� |��ȋ�~���@V:�7  W����.�,��q��e�C�jD=�Ӈ�#���<��O���G�y8��P�f�UHz����J�m�O#�`����GV9?�`��r��l�S���%�+��gP�]%����nL��1+���ef럩E������a9�S�=*�`��z�W���lj��6;#h�(��ʬtN��:g<�����d�N>�&���7�Xd�< ��*n��6?W�wqQ%�B�\o-C	Ǯr��\��IS"B~����͏{�@�TWiu|�����fѤ>����\l������>r �>���qw������?d*r��M�0 &�z�
�= ��_�����?�����.�_��W٦0<z�w?���v!���N+"�ՓJ,�Zȥ���_�ti�`�����w6U�!��P*��������P+�?ϝ��F4�~.x���!�׫��|ĴD�#Ffn-�:��h\ҟ����Gb�J��$6E��Z�{(s�ֽa����ӓ�[�)f����M��389��*�j�g�U�0���mk���&�r��I��ȃ����Seo2��/�s�%�3��^�EhN:�g�) E}I�ߌ����=�L)����A��T�0,!�p�[Ƴ\�t�"�|lSJ`�rrt���^p��8�i�:��P_�r~׻�e栨3�Iwȋ\;���^fD�9�y��DZ���g�&�Ӟ�4� �,�.#J.�)�LA7�h�u�JDޯ�9��[osi�,��ɳJ�7�i��'-z�|aL!c�rm�#7��w����o��e����6�|���:ۗ��7�N����͑�FN��zҦ��l�p��ʞ���Wa{q8{�̧9)_�}�L���6m�T�4���$,�gčy��}�G���!D�2��\���B.q�8̥���A��%�������O:[C~t�G�vZ-��!??G��ʃ��+��+���F/���2\<S�@=�/ B�:#���8��
�.��$g ��������!f.O�~t!��PB(�/��L��,�#�c����ψ���6�����E�P�3��u�}|��6�Z��w��6�O[���M�+,�f���R�iV�����J��3��o��#��m�:H6B�nz���4;�4�p�(�7��:�2)gG��g-}0ɣ���J �����:�E�k��t�w�����)>+����X�$*��T�����o 	 ��b�/$�G�H5KD9 ]գ3�"�DP�u�r���H�����k^��<�1��Ys������0*"H��� �:�!�&�O|u�����j���D"�4�G����=�ʎM%��%t���dX糎k��z��tJu�W��5�5�y��N(���5Ի@��1%���>D:�w��:��W к��j�ab :gi��Y�C:Ыy*�t��XP��f� r�Q_8.r��֙�Y�X�I��'E�(�)p�j=SWڄGbxD "?;j۬঺R���:C��ֈ=c=���
z�Db}���� *ף���VSEpA`���&���H�-�1o��)D�j!<<�P�>&%3
�?�c�^�f�t �\�$�$F :���q@���I��{�c�<�.�܍{ :����n8�8�aU��J^��u�5�k����w���K>�Q_o�ύp��z�LInO�v��B�N���9x��Q��}�c-Vǹ��YӰ<��9u�ȶ�W����������n7����ĝ��:��ݖtP�~�h��x���6����i�6H����ŧ)����9��@o�8)vC�����se{O�� )��"�.�����ԯ%��_�訿�s��`���9@ ����-�% |xR%��SH�57�I]׃���T�u��;�g&pv *"�7,s�,�C?��PW!n�Z"QR��擞�$+n(�FB���@��f#�#NW�kI�]�s_祷�QNZA� �k�K>�6�F~����W���?������[.{^��v�vX43(�#���f_�⑲	�u�s�V`TU���=��������4�^섦7�\��ն��j?��c���4�!�1˝�$9ڕ��fU�d�o�&ąiB��ݕJ��l^�[,�H��g�8��	�ȼ��M %@H B$�8 ����mn�B��5�!���Ƚ��J��7�O�*��ο�!�V��>�I��� � ,�3N����v���	�}�Ƨ	*����3�T�g"<�E*$��+���xЍ�YDT�5Ї__���(�s_���O�N?��X鵈YS��d�>�=�V0�=1���G�!�wUL�xx�st�K�^����9}u	:�'/l�j'p��3�bZ�kPT�dV�����E�z��W'�rRZ7�Q^�k�=�����SZ��Kj�K�ַ1j��/���p
���S�n�AKx�
�}�{�m�2l�� b<����W�)�x���a/�v�>�Q@�Pˠ��T�����6����,�a^Hx���,�M�@W�$D��*�#�?�ʝ{�.ͧ4���D���ѱD�%����O� ?��������1)St�>M	���T}��1� 6�$����ɔX�S/�F0ќ�J>�tp�M�F��Z���?$"�U,zR����Zo���fw�7C\����iꂙ�t���@,J�������B�9��<�͵�L�R�v��6>s��'�91��x�|��h�|�Gn��w����G�{����j�O��O�M��gs�� �k�{��t�ԔN� �w��]�	|������6�x�������?�|��/�8���IK7��/����7���������8A���7��b���Q&���`�T:!�� ���̥�Z'��=��=�]LE4w�@I>{?"	���5IC�_��5�]>ː?�>�<��q�`vXP���۴�Þ԰����h"	�u���w-���|�o��|]K:(�{Q�LŮlڳEd�N�!��g���RV� � ���i�9�O�h�ER�׷%���n鹨,��������΁ ����j�9�	��>�'���S��ȹx��`�y	����]'3&.�\6ޅWK�7ށ�~�dB�w
8ͯ{�� ��.���a.,f�j���
��ج�?�G<����!0��AY�{��,�;�E~�~�~A�B��=Ȟa����]47�4�`�;��otl=#QJ��gxԢ�����$RP�$i?o��~?+"Q^���_sұ�_Uc��G�-���?sڌfӫ}��મM������y�C��9�ƚ���p�d����l�ӽ?L����Y�ϵ�6u��r���� V;��=� �����Z��,? �8�}9�C�s�ˉ��S:��o�[T\Q�|σ�' Tp氬A+������m�plT��p� �b��7G<�	N�4��#2��)Oy�`	m<�o����Y%t��3�)�^��t�R>Iˍd|cSm��� "�������}2_Aj@�6$��E� ^�̓:�����5��k����%&���/q��x+`rm#�Y��$��t���9�V#�+�{�_	�����|�Ҵ�YW�cO�6���s�C�l��e��,\ct�f��[ך��ä���Z�D��	�d=�0���^$����I���h�P�f{U,�����J�V:����}�%���3��,4� ��~��~D�J�Ӿ��1�Q�hJI+p�H��k�f�:�el��|�G$��~θ����7p�b����͊�_Q���+�E� }p� �^��q;��`�a,H���*!�z�S�j�m�5ʁZ�@(��۾��=>T?���}mO @A@@�,�s*�j�w� ����� ?2aS�P�hޏ�'������Td~œ���9���:'�k���'l͆�,�=.rV&ěA����s�&�l�����9�	g�jgݮ��xn7�~ǁU�&�lW]�NL��Ѳ��I:���x�-�����Yw�¿�Q���?���p��4�U��km}}W�Y��QZ�\龷�M��1���t]sf6�n;q�B�Vͭ��z��V�Ni�@`"�¿�:#q�S��?���NJ�����gT|օ�gT�������N6�R�@��Lu���"lQ��Ħ�� u�k�"ݤD�6�m��?�S��=�������;�"�#vAG�����8�{���g��3���I����?�oyB �`;ɑ�y�P��qR�.��q\79n<����hC7�� XTS�s��a���@��PH���OBH���Pr�8wyFB�2�Q���j-��ȹB�TڏSo�q�4�;$�U(��k��zx�G�����!6�{J�t�z�Xi��t}�d�>���]}���IT�=��MC�:����|tC:;9�޽9]X�i����}�aY����3Bm5s���!���� �u׿�G:���cX�K:�p�o�:����q|4��|�@E$��x0(U�>���N�'�C7�	�<ٺE�^X�D��`�'ÅE�U=#�E\�?P������$=�V@d��FS�Os����y�{��'�os���"��'��׌`��<�Z �����`��N[}ڳ�6j����<�5��	��	*���;�|��K�up���Q/��9�ܜ�;4E|�@J 7G�p����TK���ks�1���+OM��HX�5I~.�LI��A�m���#)���ɭ�d��s�ۗєw�t�*8cR�j�:�Y��n?G69�Սj�z�B�ۄ�-鐠�V]W�0`]�8�gW��p5��H�A�;����9�:��F[؁��ρ����#�K'X4�J���3t-c�3�r��Փ�y�	b��D!*#��Ę��,��-������7��,n��� u��T3�{O ��_��t�ҥ���?}��"@%�Ʀ,8x����7�?z�2����C'�Pw�zz:�C�a�CGl�Li�	u}i_+]Pߧ^�{7��=���^���B�Z���'���R�C{I�cH�R�Jm���،�kA�\��ݚ ` ޴�ta����V=j-���?d����y��u�&ո��3��DI6Q�^��_l��m�&O��r�YDܶ'~aD:Im���'�ߨ�r�.s�q��}��vo[9�������B�2�����ap�Э3f,}�0�!|��a�� SH �����4@&�"�;�>�h�~�;8p��ޡ�9z|�f+6�a�C���} z|�[A�c�=���:�^������Z;��#Ѡ�H���}�|�[	!�c�I��T�K�x�eT殹�$Z#��Sˉ�%��)M�o�@��oJ7�PTP��m�c���H����x7��&LǰǠ4%>��H�t���3�B|��W��zP�4�os�<9�wO��nR�j�̳�M��� ?N�I[&~�㏸{�'�-�W��pV�V���(�E4'��g��zD�N> �A×=L��i`�f.� ��|�k_k`
W�P�@�+�.�ؒh�x�������p,s�J�'���^���m��t�M�+��+�;��{��Fd�)� �,}�,�Z�|���(�o���5���˗/���P;1\"��]h3Ok�<�]GiB�/%/ّ3�=o!���\�A$�*8���|�g���!�P#�^��V�ބ��W]yxv1�SUM׃�IeQ9�;T��.TƖn�q���	@`�o�y����m�q���nu�|�|���+����.MN��/6��:�#CN���ր��T�zG>�~I���Z����� ����$B�,V�x��'Z��, 2�a3?c���,{���˿�KM > ��:@��`zI}:ʢ�^�����4��� 4�H}�;ޑ^��a,��g<��²j�g�_�	�F���}�g&����]�#��t�{���!�ރ�>���nP5=�я���bE�H���灑�n��z�������>˾��\�pD�����!b\�R{5��U��{��?Yo�^���_��4�NdX�iP��3	�}�3�n}b�R��\��-�>.��~�]�~W�u�o�F'W���A_'?��Q��~p�8%פ4щ�t����(m�u`�;�ND1&K*�=�7m/R?�[��I�2���%���?�o��c��Ur�P�@��hV��[�e�� ��8|H0�D�Z�ı(������A?��TA p���&16u�7`���g7�����d-�,����t����%�>��D �>���Qw�	<���� sH0	E;@H���@����H���׈{�5v��J�^j%�7ZU:��<�b��5�Z������1x�3����Ų7*��TZ{�'�M���}�Բ�e�8*����YG4N:\��r��͸'XW��k�:�����~?�or��'�8���4�;��������1Іr~J7-=���L���9� �5?��Ӑ���3���,K"��oDxJ�Ʈ�x�A9I�ߗW*s���s �سpÀx�����#l!8j,x4@��0�*D�z�3�i�JK��4I�oA�u�`G��0�* ��P�Pώw��3V/�	�CDSPp�(�� ��F� 6h�Q�8�<�r�*1�;��$�Ɔ}��i�>�'uۺe�`zI�s�
ƞPx� 쉋���$73���IJU�ޱ�u���a�3�
�mky���r�R�{_`~l�o��a�"4rVd�7�j�����0��o#i���|��W���dtV��7s+p#�l���uץ�բ{�,�+�t�n�Q,ĉO�c��ޒA'���^�ȅՁϨ�E�S�醟�/�"�-�sX�=��!.uUO��ԟA�?�.�qx	� 0���wC�CK�W �t�  H�-7|��}p�� y��&��y�q��C�_sA��N����xe�E�Y�3 H���yQ� ���*���gji��&�Q%�qSO�sB���R�e?�U2ae�U���~�F�K��Щ�c�c�y�Ŷ�!Ǆ�4Y�����B����^�X����,on�<��y���m�A!����n�6qc!e���^�w���:(�{��^�W#ߖtpN_�;y���ͩ���pB��z+�HS���-�����[�q"*��Q�H��RD,|^�T�ċ��]�ࣾ,�����^$z���OA�t���i}��eS����]9 �AH ��G�z�?�`c�O=\4x� �[䢹)K���E�Z�����G��"D����Y?$�'ڋ:��T������K�[R[x"�DB�Es�K�q����$��ҵR�Ur��K�������wӰ��!�p�m���L�t�O_�AB��ܙq�g ���#�dS�]�&�A���D��%qij���ڶX�gy���z�ʑ�� ��]z<�n�:�<���4���6������K���}?���z��1-�4m��wT"�ఈ�\2T+ }��e��?�0 :�<t�FSO
|���V�
��@��kȗj&F��w���WF�ȓ��zP7nF3�!����N䢹P"�~<�=?�"� b�\�2Q=J'ʿԆR9��oיW�Fks���Y�d�=�˷ga�X;=�iu��M��k���0n���0Ŵc달�H�$bE��BB�d�����)T��4�N�jeR�C���#%�@O�Y+�Ivd���S���T����[�[*:��0#О�]����s�y-�t����l�"�׽M�1��w���/�]p��#1l �Q �MB��3����A�� [r�ܠ�*�\�����<m������u�'�K<)�!�����#�KՓ��"���{iL�6ڑԥAā{n>*[G㹋i)����X��᧗��މ�i�>Ś�{�R��#g�]L���e�+���g��kG��K2��k\k:(���9������&������H4=�mz�_�]���;��|�S��Á
P��`ڠ,��:�:8�q��qs?zG�E�~n���9�T�3^�T3�+ ��v��רr��$ /� ���w���5��A ��A�z׻,f����C5��~��)�o��o��`�	W88E��\>����M?��`���p���L���R���,���G�s�9ž��G	���P��kl��#�r��������~3���=3O�b8ܫ��^��������_���|���Ϫ������xu�b��j�i��1˒�`���b���|��#\�_�G�8|�<5)��D����jBX(�?�����&�W���ę�'mM����ϫ$O8�7��̥�8�}����F��r0�I�F�y,k10:��iBI@�����:|��&6������p��!y�`)t�����|ի^ef� 0�J��܇d �F?��?jy ��v��
��?��`�V=����͎��'J4�G����
p�D�������nss�yD�K��%	D�fԖ�s��j^�-r��i���=����T�MSV���T�=���)�z,��]<%�s�}��@���}J[��+':�R�fE�`��Щ f ￣���~�����jT�(�¤�"�v�D��%1�si�|$xND�����ā{k����-���(�������'�s&=���=��i1C��OF���cHĿ����W0�A~������q�|����/_��.]�du�A*��Eǉ�(�� ml:�u2ʀM>|����`��g P���(i_zis���u��:�J�D<�i����ys\J�����������.�f��:��O-����Y��1��
&�A��f`��Zan��?{,�����뺞�&�o���i�$���t�$RA��o��Y�k�k�Zj1��>�r����z�~^��r��,�t~�y�~�.����$�vڗA��R~v�M�2�:�O�J���$�~�b�@���KJ�8�(jIA<��MQ^�'6b��O~��lp��v�8t{|H j�?��U�n�8�`�_h�p��Y�e�^8Ջh\��2 I�"b����}>�� �%І?��?H�~��-\#�]>���A��#��7��"p��һ��9���������{���X�ѫ~�>L`��&�w(��^N���b�����q�u���-z��0,��O`��% �[�~��`���{j{���VZ�G�����������t�Q���U�u�]�d?Ӗ�Yg�܌6=��t�{��1�+l��ӴFlʓ�)�a:u�|elzε��+h�Q�N�Ӵh������_I��?S��d�1���8Sg�xoy��*mF[l5��gHDҶ���2�ɟX���H�o�W�MF���"�:h�t�y�X5c��Iۡ��D��ڃ�I5�nfњ��~:D��8ip� ep�P��=�b�t�C�7s��['a "a�S�@~l��{8m��w�3��>��<AX��� �
��#O�H��\���5չU��=��<��':��(=���,�P�~�J��d�i;u=�nt�&��D����#����"��N�� .�q�]�����#���-�ܚpp�H'��\\蘈������U�p�>�\�	�N��M��>�r���6�t�W��7t�\�2�����9;?�>��=��M�6����dj&�<a  �Zg�M�H7�	���7����L�,+��C�i7w�eF���V��F���4U��}�9Y����-z@�BZ�T"��/\�~֋V>����%}�������.eBr�3��7�a�z�t�Iؘ�t�Dk!<�����<���5�@@-����l�{iy2Q��O�J�Ӄ�A��7G�yz�4��X��W�"-S�`�,_7/�]���V���!���zȭ���vv2)D�m����6o�u^頠v=�ӻ�Y�~�������,�9��hx��ؔ�7���
�pCݽ9g��Z�Z��K4@~����=iK���l���H��왵�R�"p��3�Q��jC�}�]��\�E`။�~��`���k<y�86w)) tq*�[�d��>��C&L.��DV?��� H��{�[�bV=�3 ��!@����o�;|"#���s(	��r"�h��K�>W"��9��R�J)Z7�;��R&'z&ʿxF���@����̰�7�<�*�t6���x���;kз<���1��ufD��,6�䤦��"��Í�g��`���d(K��F\A�D��F�.�\F~��<��ę�:��2�o����d.���Q��D�H%(�#�6�`T���4�ϬCҎ����� ���i/OW���5�5���S�������s�رG nu`HF���:��>� p��.P7��>$J´BbxŹ1��گ:W��'�X��K��#��E�}ު�ѹ��G�^����:i[�7݈y@�zս'�f=Q3��G�ߕ�i�K�BP��w���>����H�%��^?[zv��Y^\دx��؏�2�XX�m;t�cg��d`�6P�E�G�z�H~PJ�(�h�2�?�g���kzo�Ő'[|��]�W��.���6x��u���* .�p<�Zp�������3k�-L3��ۿ� ����������M�Ka ���IN��J��M��eD.\�&5�zA@���9*�0*���{�T�������w�T�7���3�Kc��)ͣ]�k�$10r���l��m�}>wz����1٘�bY��Y�
�����i�+9Bꙿ�L}��D;x��S�Ǯ�H�=�6A�%խ�*?�z��].�5��<K��`�l�u���R9�N�W����.�]������z뽨�R=|;�\��{Q��>�! }�/@��= Vp�|`�[$8X�-�78���0+pݰ�A��C6���.t����}H ��a���]����>�?����٣n�	�?Pa� �9�ƹXJx#@�c��zݿ��Q���њFߟ��W�ѷ-j�\=�&��?��˒��u��E���d�1q0�?1�հ�Ԅ���<�tX�61�[Mg�Y��f�z��i�.����$v'��_�N�^y@z���_g���xTSP���Z��e�e�;�s���l��~���.&���,K��W�e̵/�;���Ԣgx���y�V<�#��_��_��雾�@��o4. ���˗�d���5T8x�*p� v�i�;�{ >�8y�������ນ�4+�$��[ }�˳
���[��'���g#�3�K/A���3<��#���1�:�K�Ṕ��Sߋ����홫���{�Jp���?5��)���������y���؀��o79�n�*F&td�Q�sT觏��5���8���M�T���?���ͻud�	f� ����z�2���k�'~�D:�h2�*��K�8�򉸙�>��#(�ګ�i="�(��2�~־�B�ǖ^/1��YC?N�K�� ���@5#m�c���?��;� ְ���_�U;i ǉ\p�8��>6���T	!C>x�n��=�w�S�o��A#iy;?
�:�=�u^\������i�=�_;��s��%�m����=/i�IK3�a�40F^u�������=�Sy�頠��-i�9I��[mo]ӵ#���tB�9U5 =�:0mG���30`p�����yv��9��kP?�6�8B�q��EǕ�������=zۖ9&ϵ�$ZzUMdq�����b�orR�Xƶ>��X��5o+�D�k猔��Ķx�m-O���YS	�/G%�K��r�|��a�]� �� ���'��=�� * P��>#;�y�}�`,���)�1��A,�UH�F��sd��q�3:���ύ�a�`�@���q���Dc���7�� �9^��uM1_M�7�x��7��ո�M"3�B�����[�:�W�,�Gf�����{��s���j�0+��Qo~>�ƨ���=J���3}L\+#���y` V}����4�Q�lq�и�3(fk�ɮw����@xs6�PjG�S�\h$�J~A�w�����%�'�*x��EĠ���%.1���~QXm+��`AGkx��>��r霍\4������|{�~�4��j <��b���������: 6uQ.�Cp��<���a��}�ӿ>y��c��wi/�0K\�2,O�7JQ�Z�9�P˜�_	��׮����&��/Y4f���Z%��\^�&�%5[��=I[�n��\��8D��b��Ů�G�/�b����c�f�ڳ�0 ����m��j�Ǝ�N9�^�S)y���H��K����ܘ/�o�Ee��3���d�$�h'�_�*�hk��ZM�Jc��R �d03�&���N������J��q�y��Y&��{�^�.�������{䋼P�E�ƅ?-wh>�w3@���_:V����%����֗U)-�DL����h�2y����0�a�@c��,�fa�__�J�./���l֧',ð����L���Z��c�Ȼ��g:�ɦp-�o@6c�3i�,x#��lÖ���l���")�9�y���?��<�x(ږ_�>������ك9	'�G�ݒ�S�&��9�P�G��Dj\Á)�ȅ35p� W�G2�
�5�p���,G�H<�K_,�������,���C}��4�(P*`;5j�?���K�/_]?���Qb4�-���З����/D]7^"��R����V�T\s�_�oN��.cr���v9���) hY�����mI�~o%�,�Aå�R�˗S���+loΪ� <\��)c=�Xu 1��)1�y�.�+־T��Gѓ���I�&l0���"~\H������R��ez	ƃ�O~a�u��LΜ� �pn�����/7�t�q�����g?�i����x�9d�E���|��������'�+%	�M�s��/�q��������,��y�{�c'ta)t�ҥ��W�������A��+���۫�C��O%�轹���fn�T�T��=s���>in^�I���LgE�XjJ�Z��g��[k�o�I���\,g���L��������"l[���L}nB��\4��&�G5�A͢{5�Zo�zcP�T�XX�:}��	�>WW������9�X��嗬4���;���K�Uzv�������x�9��DA¨A����3&N�\�	�8p��w�� r��G��=V�yx�|�k_k ��i�r����~�g~�|���<�9�K��KsQUW��OK��(�q��/�Twq�ڷ��9-˯��P���ќ)��>y����󌡹\E۫p�����~IjRmD�9��}�Ib�����tP�W��8�Ӄ�dtd��r�i�N�9�h���gk��S��z��1noQ���eK�H�4}��ц.�&,'�ݮ�e�I�'�U/_ר\�V��x5�>��G���/j�o;ǑB�O�5T)�kЇu�-���,<o2�g>�Ƶc#����,��YW�R�jy?��O5��u :ʅ����@�x�Ӟ��q�{�?�1�1<$,�?���]���~ÐDPAm�!��|�z˙hL4�b`�����-��K2sR����Y.�D���l��m���H�+ک��z�i�ѕ�P%���eɬ$���Y���wB�ӗ���H3�o�c�G!v�����E�z��}�L�@����i�g��y#�
G'�_|�={�y�K,mGm��������r�%��s���J��\��d���5$��s��K�|�3����/�������'�������e��APC���O��O��F.l���F8q�W�L"�����2��^��!A<pu�Ր��y���j{���+��槎ӵp��Y?�C4��<�u�߯�(��/�<�ǜj�xֹۻ}���Sp��^bS���5�����ʏO���頠ay��n.���ȼ]����i'/S�����;%���KS� ����uլm Z�M/���7Y�T�b��O�ujWݠl��Դ騾�E��u]��Gsԛ�j���OG�uZ��]�:)�:3QC�7s�~����وm86v����Y�{��n3sY�ƸI2޹��綛`]j����C$�)����_<["�Mk������(�� �}>�^ʍ��&�� �t4����r��U{t\G@�N�8����x����G�����CE�kp��Ї>��9H�L��� ��>���s��MdZ��L�9��9p��0!���0�Ļjɥ�5Ε��8�B<�������8ݾ�y����oй�%J%
:��<H�Ą�v�1�P�����3��ז�c��tښ.!ٮ,�y���}?���0�cVq����ͼ���eu]����^�<��C��tK��y$��j�W?��vy�)�6w�^ 69�R�U�&-Oa־�� W;�b�.�qX9ކtX��i{�2)�ܢdm������Y�Z�ΛlG�H�O�?����I#�B��'�I�9�d�vɽ�Ý~���Ҥ/ձ�{N��'�S" k����{P�4�n_������3�N ����T�K�?��7��V�2������E,�'>������ &`N�>t�p� w� 8<@F�K�[�j�ԉD���p.��R���辰�8�}�KU���KǊ�鼧̫$xm��ʗYZc>�5O`�3s{fVϙ��Z������)�;.#ij��(�i��oT����>�G�����kuY�x�^h��s��L
�kͼ
�����naޚ6kX��rQ[�y��N�Z�mmt�΃�n�zx~⫪J&����}�.~��!'VqK���h)щ����E�<s�S�������R�����>q���U��� �����ַѡ��;   X� _p����e!�����ߧ�>���F1M6Q��g�ˇO�:��~�˛��f��t��kt�@N�R�&�9WJc����}�@9�OJ��K��z4J�"P���H*q��}>�|���lq��<p�`
��2#��[�>��X��:����Y�֮!�;���i��t��l�������	�gj7�NN'��	[ȷnৼ1OO̧�`�XJ0���֦���ąM��}
`%�~�I;�k�X��oGT֮���ХT"zQ;|���n,S�����[Z�0
��K��K�f���"�����A�����f�.� ��%@�<�S-���`�p�H��Q'	��R~���G�� |��3��]�͍R_G��K�>���6Ǒ�#m���s��KeD�ZDdJ`��?���;3&�6�з��De�O<!���5��5c֮tP��Ͷ*��@��`	W��}Qd5.��Uo����3��]���{"W�7mo�|���b?���[�g�����������G�܏�G��[4��%�KS"\�E4G�JH��J&��xi�5�;��b�5��8���y* -t� e�~��_o~��?��4�$"A����� E� rs	栗/_6���x�R�
�������cD�xJy�l�����h�UA���9�;�~�{��}2]>^E�I���#��?�_:7������B>����v}6i���M2���ڄ�=1��f���ׁ��[;l��I'��Q�{�S՘O�Ox�g:��a Ԋf��� ��g�=t$s�(u��y��]3HB�2(p�~B�z�-O'|��R}O����`Z��ͩ��.�9�gN:�o���E��縬��<&߷��\:�r 3�-`��t�@��*}��y�5��ì�xz����	�������4X� �1Ku �Moz�9S���!u��f��Q_x�$��07�����	[������c�[�ϝ('Q�f��S�sܺ/7���*q��P�����a.��D�l�k:e S�-�jiW*�����\K:�z�Ik���s�2���/�C�_w�|k���X�Z]�f�59�5&�Y� ���ą�7�p���v%?Q���A�YϾ��W�D^��܋�&H)��$-qb�s��c3mS��#�\�^�~o'ϗ����^��}<�x�Ǥ���� �t����*�����0[zp��" k��`B	 �Sw����tπ�<�я�{ p���j
'|A0�|�;ۻ�����Y����=Z"�3'���A܏�g��F�b�����*>W���w����ވ������a-�Q��������~:K��4{
������ l�:<��hϺ<N{���X�a�H?�����t���5��`@Y/;�̖:���E�������w8(����)p����Da�e���Ʈ���J)\��fRjº�]����%
___�ҳ�W:cP�F�5�N�}p�^�����m�D�zғ��^�������8����1��0ޥ��C� |3�7v���s���0�xz|DԺ׽�eC�4F}`�˿��f�ύd��G�]���IL��Ѥ���j��h��qў�O�H
x�a��N��<c��y{�T����c�OJ׋�0� z�;IZ��|��F��K}0=�2j@n��O�I}�#es)�~G[��,TFa.ެ{�ڎ���V�f�v� �����?������T@WN��j�O��e�`N�J��X������M�Z�ͭo=�AZlo����1�o��#$���ͅ����W�"��kg��Qr���z������K5e�4����K�ā~��p�T��>N�ҧ˥}>�5�,�@�v�7��lHo�ۍx H ��a!P�:{�� �!WO E������uiܙ�J��̇J���c��N�N%�1�(���
�y��u�7bvx��u�=��<��T�L�
��@��Cg�콶v��j��޽�a	�C��+g���E
J��UjR�ev6)}��Io�'s�<�q^頠��9�	�ꡐR&;8r,n�4Np�ߢ? r���4�����C�{���8��ŝO�x����b��iG��sȑk�hi��>���$	����9g��OD�I���{N	�J"0F��	s��q58$�Z��Ǎ{8(EGjT�9�� �:����>�-���D摏|�@�x�.j���K%�HZ�>������9��y�5/F�Z�/?�ڿSItZ��!�+ZJ�I����ˤ�$�D���HNV��i "����lU��t�Ҿ�cb���';2{�~�9�z{���lx�[ڣ�jZ�,tT؄L▜����c��ކD����E�ؑ�ܶ��bӅ�4�S���sC�J�%�wn�x��sqQ�ʱ���K	>$�N�(�G�a�b����� ��C�߹Y�g��a�-ܧGM|X�Y���}=�<@	� �������_�Ŷ B@���OM+x��hZ����㹏-��Cˌ�Ń>���噌R~���Q���84_%~�M�nc��ٜv�<�*���k�ҋ�E�4 w�a��-����!Z��V������3tBu�����ȝG:�N�4X��
���J �E!�`��z�E�Bd���u���-B3ʞ���s�0Ej=��Ij��jk!���j�z���%n���G\��|�����W��J?�t������r䌀��
���c�bs����
�XS�����6y�<�2 x� Cփ���*���7#s1 
�$p����}�*i��ٷzͻ^昰�"՟���:�DJ����u����W	Į���U�V)&�gC_�/+ɯ��iZ�ն�aN�UM�4�m�k3����?x��ݓ���Mnh4�;����o?p�����E\ؽ���|�����:�|K��i:��26���B�j�8(s�.ZN�h�����r��m����@�W�(��wT��ū J`U*�s�� ���`#W�:@�k����8}��|�q�x\6\3 ����7L�����x��k��=�9����|���Okԏ��x�qy���s ���ט�3�t�G��y�~�$�9F��K�ۧ}淖�K�  �"IDAT�9���8ĥ��ZV&�*1�m��/��n�kO������ �ᛎ��a6͗O���h�6FՖcm��p�	�>Ć��#gE����s��r�~�]=�: 4-Y�׉uU͇��#���]�ۿ������DGb��Q*�΀�|�d������d(qMz����3��!�q����+��S0�I99n�r��`�����]z�_�����X�<�Y�2o�඿��1=�y�K�x�#���=80wˌrōc�?�.���3t��ks����Ãw5vo�������g(�ߕ�G*<_?'�ӗ��#�N����\TV$D�#������o�͟��q�~�2�_"4|��T0n�����7}���
�I}��I��� �U���-o��o�ka/�����;	~���bAT�~�8�8�L�1���>4
����怳�ʑ�8}����ไ(O������S�%�pNZ(q�\@����8D}?"�
z y�'-m�U�a�@�p�v�7{pm�
�;�{��V�هM?ʢՍnjj�b�т���V��O��YZх����u� �}2��XE ������I��qQ"�	��U�yF,�F"��C�|F%M穽C�:��p���l�t b���"��A�8���rc~��\�-?��G���6��	���]�>@IgiW?wBc������7��1�5��:gm֧e�,�zz���9ج������4Z�>@�:�ܬ��k�d��xO���\J$���Ӆ<�p���>߶S@���h3V����k�U��3T�P���4 �k��k�6 v����x ��/_L5�O����ǁ-�c���R]�>U)`O�i	�9��\G��,�}�}�MCӨ�戳�g$��U7Z�'&�a�{�@h>��{%դ�/���j�S��Jң?qoׅQS��g*ž�6�����w:�?��K�1�:� ��������ծQGiY_���c����G���Y�`6�u{�#��r�PK����韮s����4���Et�T��KYۤ쳧Z]5��Zu\���  �nޟ��ߕW����D��j��$"���u��׉����aB�Ӹ��"8&G���<���L�v<��=O&5�,k�6�p��	��,��U��Z���A�;������K]e׳J��9e�ˤ_-��,�z ��\�}'������Bǈ�D�9��"<��>�������#���.����Ӌ^�+����O���L*@{0ӎ����7����E��K��)η^�2�HV�����M�����N�n�4� =Ǣ�f��E M)9�5J���w��L<;��<P����߀��#M%P��fG:2�����#R^��8W�4�˰�i9>(�'�J��y�͹nNuK��n��[�3X�-�ts��#`�?:.�����"׻9�ة��Ҫú���c��������t������T�0���q����$��2��X�W��t���t�����_���p:�tX��}�3�T�ʻݭ<��'�4nnQ�#��N��j���� �o�4��J��(]W�����kIZ)�m�|����X*cW��I�������e΍A�^k6î�D��zP.��K_��!����]�x�����t���']�ti�|�i��	�^
��ysT��m��>y`�
�*��^��z�o߹�k�瓗�	�S�Ю���qۥ�����)rb��L�y�M��N�F�3b�,@�%�|� o�HԮۚ��� L��Lx�D��f�a�=���ˈ$�]����5#���;䛵q�J���c�-Ҷ���`J1���>��X?��@N�]AL�SiQ�Ri�F��ԧ����{JE���*����RR��mr"^��3��G���E�گ{����4τ?��E��*���W���p�a��M�8j*��C�&�~~F���?�u�6-7꛹��O�����.�����T���4y��R*��y���v�C�[,V�2��Fum.o�Z�2M���Mv�h�T9��7ۑ��+�s>���'�3�yJ)���0Il���]?��A�.��i>PU�͕���PN� �S���Hj�l	XKz@}O7a���|K�>�r�z&��1GhJ����j�R�F�� X��g� �����p�n����t�ЇG�Ͼ�݌��>�ˇ��#�%���ID���|_F����w|Y>����)z��+j/��L&���������F��qTONR�ǘ,�M}o�<Ӟ0(��6rO�4��_nk:�����>�\��-�Ӥ���KCA
؜u���ǧ����yfe;�ŵ;�"�o���M������s�<�G@��?A9�,@E�z7�S��~q�:�a�J�����V%��J�e	�x>�� G�s�0p��up�pu��?��ַ0ͤ]?OѢ�p� kx�D��O���6�[�=�������]��DW���~ex]��d�Y�ߨ}�w4n~ND��~�U~�Z���:~F�J��a�M�Һf��qU�����Eߧ����%�Ro<�O�c?뚉�`l�h��y��;\�H��]�ʃ5��3JYe �f{B��h��G��FU	s�_��Q��h�G�)ߏ�3�Ƀni����i	 [�["Z���6)��3�#N6��/�v�K�f0�W�����=�Qv�Ox��ͷ�b�>�� r ��_�j����x��n��#F pj���'��~���y�g��n$MF�ʐ�͏7��[���Ծ(�	V\c�Y}����vd�8߬oO�TR_ocӎ@�j�x��t�g�30�i�}�X�p:�tP���̾oڪ?����Z��4&e[L�&�k϶�����땮?a�i`��Y�*�6������3�q1ԋl�����M��[� ��G��@?+�:�N9io
�ϗ�\Y���U��
6��h&�T\��N�K4Z�]18O,�����S�N�17@��*�>8y�aF�oѸ�M<|�n^��q*����nRj_�q�c4�]��&�~lY�/�ϳh��x��8)+M�x�J�i�N��{)��MV���d�ӊ+dn�Sh��Y�F����,!�Y� 7m��l����
���)g�,V�t�m�� $��<��g��SQv�uz��O8�v��yO�9Q�@�����=���i��.��ӎ�s�����S��G�����D�}s���p#W2�����8��xe��1���A�y,y
�����?��?3��>:x�=~��8�����'�����.�[��[��@# ��{rz�%��=�ÏO�Խ0�G�}{#@,Iw��W�̩'�JG�������Ku��S4>$��[�][�D�ٷuN���Z^i����{f����u�׺zM���*�����s�]*3����TՃ����>N$��n������m�znN��F�,m�'�԰���y̬z;uv���:�Y��xu�o���v��y/ ��0o��A�k1�jbp�`�s8���:X���CT��m��}?��϶=��`l�0#+%�����;m����<��"� 1jc&�#'�qg�)��E@��<�)v��}���v�
�����e�o}�]ů�������s�x�����k.��~ԋAM�fH��Q `��׿����j��YU9��c�|	����1*M��2u�rXO�b����D�������="������? ���~���Y���z�{�`�7��ۡ��I�ͧqi嵩ǳ XG���n.�7W���z_U��O�����D��`��3�IZ,}��Y,BqvvR\��%ܵ�NZ/������_���G@�X�4��}����I�l�-,K�FN0�x���iڨ�K��o��KD���K`=�Ex]˚��^#p �0��}�,��O�}�k\��e�UT=H��n�����$P��a;�m��q�o~�x���_$h��p�,�s��{^U�<�9���O*��&�,h��0�~� �|�Qh����'�#��?�ʥ�S�τm⽶�X�!q�I��Eٺ����6�a�9��&���'�R�k_�]k�z�*SP\���6�g����W�;�!���Gu�C�mֵ=�͞� #��8y���?P�U�@�s���ӾC�Z��>�"8���U�K��/�/Bs�_j�\��z]�xQ�t����w|GVҕL5���u�}o��6h���� ��@�D.޳E:D�*�uW��0��,=G`���:{�D_�Ҝ*��}RTy-7b�T2Rf����x�j�-���"e�`���~Yv��90cﰻ���R_���$��4s�u�3�ՠ������ؽ���w��3����pڶ�v6�V8���i��E�߿gT��UGdV���%��m���x.�t�D4"�DOU�deڇ��vxnG��u҅Z� �|*\hsD%�X"s�AX�o{�q\��!k�]ʑ��MљZ���A$�Y!�|���c�4AN���oG4O��=[�䈨O�)Ij����/�OT��ۧ��Gsŷ]�9�)��MĨMޯ���j!iM��iĀ�-��b]TB_.�
����F����7�א���w:�?�� ��j@a~�gb�U�˷]pPʶ|s��6��a����Po/�����p�^�тڵ���+-��_ԥ�yɛ�i��#�����#����qI�0�����g��J����an	���qn �h3����t'�����u�����������+N)[h�>�<�{��o3UV���"`����(�{��2^k���l׮kM$�`��*eF���Z���3>���_��E�1����z�6��J��92l���������?][��'	�@L�`��PM���n���l�d5�V�G;Z��m
y�d�$n�.#%(z���']ĹG�e�QGܚ�����E��)Zо�Q~l?�-:B�,��虨�Jy��"#`��� ���h�����Y�@�s�M7�/��/��������Mo~��=�������`�^ ��#�!t�������)]��O�0P�KN�$��zG����	�'������]`Zbh|�4�����9mî91S����A��\P����$�z`�����bu��4%ft�8���|Ni{��ޯ�A�_bHok:���6w҉-����: )۷���A���6vh�������e�1#�b�|T���r��O�ҁ�Vw���h�� ^�G�XI��`��Ri�Du�q%0�~��>��8m���_��W�/��/K�w��o��o�����L�y�kҿ���[�,T����f>y@ DD��Ozz���m� ~z>�>�,��i� �?�ݗK�\'���=1��K�P�&�t���LA�y)�?�/`E}��_3j2��?|�Q+q�ROtVO�-�����	.�i�a�K� :z�����Z�M���5ͭ}����wmG��Ao�F{�-�/w��wH�Q"��^��^jb:Z�����s����M:���}8G]t�w�8�ۚ�MEyF�%~?��'���*���C7�P�<��0�Mp�������r����?��f�kl������!��{8��΃������w�6��8|e<Q��
�sDZ���F��慪C��'6��������+���C���>�p��Lu��U�^]�u���3YkЁ������?9Y��:Jy��:��$���w&2�M>�0}�=��|R�4W�����>[����F�6�OH��Q�T�>���ɇ ���D��S�����t%����Y��[xm��y@��3�Bsd�.O�C煓�`Cus�x��i]�u�u'H��4�ښ�C�Ӈ��7��D���T�4T�L'm�KGG�@�C@H�&�E2���� �H��Ci�$s��Ѽ"��3�ؼ���q�.U��ih���P�#��s�mE�Z9����AZ-��������/��S����w��g�{��>�mo{[��xw����ށ�������t������H�K�G|��};�Ѥ�Toիy6���Xۢc��{o)��N�ϛ$r\t���	��楼�@�A��(s��ı�m�3_�7�70dU?�W��q͚ �Ő�9�g�od_P��'/��'k���%�z�I'��@,ۮ�[������{S�����M>�a�ճ�iYe��g�c+���s\���t����[W���OJ�w�P��1����뺹���GU�['��6���bjI܅�H}PBo_�T��;�L05�D2L��HM��0P�ؒ��Ÿ�yN�9�/�R�����u�״~Վ1�t������@�xS@���}�ķ+�y. �6� n���ؼ��/��\�q ������6����:��#Sˈ���?�V�cs����4��I\�;����4W�����h�;/�h��1P͹Ф)��R	�G����FF���=/Ğs�<�AAi����7��i�Խ�����p�9�>&�'�~82-	&��=l����ϗ@S�+Z�ܹ���ݏ�{b1���<�����?�Օ�� ��r�s��f�v�L=iM��.�_���F.���2����,����ri�Ńa�A���Л�j9�[ׇgV�}�.1����G�z�8E��Z�`\"sI����O��e�%��3��Q��Ɉ�Y)69*�ݪS���2G	f"u��Qܪt��u�r�v�<�����;}��I�,ʝZ��iѼ �I?f953,�<	�%�}��<����]�..j"p-=-j���:�����Ѧo���'&��_����$^Ё88�O���d����L/y�KL����߸3�B/n�)AT�Pd�T�R�u����s�����C�J��"����y_f�oᙳRt3_^��E��jG���T�<�=.��Կ4OHpNO�tz���&��`g��Y���9+}�d��ΝXo�M��T9`��-��؀���~�2b�4��q�>i���x�O�]R�1�%�����Nv���Fd��Or�z}+�ztcP�C���k�:2qႻg<Q�P���/��/v�D ϙj'���:r����� �~��ȿS��|����?��Q�s��^��P�����_�R�D��笮M�Y���q�%�q��p����l���f�m��¸N�ڑk����{{�XP����&�u�\9���Z��u�~��F=�q푔s4 �u��2b|ʔ��Ջ�Ly�l; ����	�]M��x�I�O^�8�'k���2&4��~��}�Iy���;�y�Z辎:>s��փ�T5\Ȱٿ|�rz�Ӟfnh���ES��R�{�Xz�To��&�w�/�Mԧ>��n�|v�]u���Kg�ފ���*��f��i����$��{f�@��{�M���]�a!|�����I�𳏝��9�}�->9yg���Ic>�OV25�~�uZo�9i�;�'���W��V�
ދ��(�s���ҽ�Z4�#p.�h��TR�(�yN��*�S@�m�4x;Lٔ�^_�Ј��t���o�fv���y����G�|��8��r��jK�
�^d��s��O�����A0� �{s\��G��ޟ#F�	󮗽5����R���1J�z;0�n�f)����h���2��f� �q[�::����[X�|F�����=[TfѶ��IW��WN�g��I�5�T�h��{���dJ}+�<CF����џ�@	�ǲʢm\�X����r���ō�8�Ht�7������d������?[�� I��a�w<�j?� 6d��'�y�xJ�-�{��^+π�^��fظU��$ڿ��h��}q�:f�}�`?��Ʋ�K�2���:�J������֟}�g����U��h��kAzW��T0������/��~�L�K]ǆ��0��W��~�ݿ�\����;]�V��ٺIGU[7�A��X��(_@�I�`�����A��+��,��������:�U?a0q��=뤅�䰆''	���?r�5�������乸����rO9A�W"B���P	�r�~a�(d`�G̓�0�oJa�j}�<]��3�9�r�ؘ5��:;JC t�ԇ>��o����5����-�-���4���?��v�>ө�'8�4�������J ��I$�S�/�}�ӏ��n��� 9 X@P���u�\��#si'{ ����V3?#q�ۮ�6X������^��MI�y��d�1�߾���s�w��1@��W� `}�qk�Kf�ts��gr�:�
�7�A��=����������v�|��W��sJ����}�:��Zބ�'��3�N�E�y^?�|2�L��wJ�ț.H$�MyPb����P@�tP�ٕ<���c�JRD�E���ߧ�|.�|}[��c�;��[|b� �Ʃ[��}��o��/|��]@��W�����_��u�{]z��g�v�4�D��}���#�N��9p�%n�&��|�����S��N����?I!�>��R?�6��o�.)�ԗZ�*�6M�í浴�C}�O�5zd5F�]LƄ8�Y�s����>��+X���1��M�4�����E�����M��U4K�W	�Xժs%G�u�[�JD������6�G'K�tnA*7q�%�w%.L��w��Q�"1�\�b���nz�$i(�i�h�_}&�RIn�t ����#!`�g�g�w��a��|���fX`�M~3J:�����s��n�?�疀1�|4yЏ��`�y�JN�3�9�$�_���Y�h~�6������o^�T���;P��0USlX.r���i��`�Ǔ]���Y>��n��v��Æ�y"�-�w�q����._=��J�+}���3mQ� e"0~op���sS�׫�����|3��4�g��35�X��i�!��6J^s��+(��_����v�t�~����kN˷÷U�/I<�(�S�Їz��>���]�z�!��c�Xs� u�}��e�߹���m�~,,.f�i�X!Jp��_XWUe�\��b߱���+���c;ء���q�m�9�ut]��\	$����ښ����Q擿M��]����$�^6g�?6�����i��	� g��x�v2���ԫ�o'��+�{�4k��6�yP4�R��q�C�ُu��mv��A��N��Hy�e�ui�v��i��A���S}R}�� ߍ,����uHK��x-���*"�H�������!�	�X4��Ġ��u���o��]-�ϥ9bq�Ѧx���R�k0����}ޞ������O	��\�0���|Ol�����w��QSM��vm��k5��9��yn��M��ڍ�}0���f�m> #�+,��n�uewLǦ������^)}Lg�4] ����� �uf�������8X�i���@��y��ԋ���{nE�@�y�c�&y��K��\��z�XDT���)Z ��x����>�r=�`�����W�qC��(<��1�ޟ�F\�0��{��i��j^�Nú�%�%���w����%�h~i��P�.j���h�(.Ϳ(�����i�ֻD@����&w�}��s��Z��o}:lV��ŶZ�~�/�v�/3�c��s����n���c�{g�����t�2���N^�7�{��0��xQP'gVe=>���E\�<�u�ܝ�'��J����d�<�Q���o�=���;�["p,=��F�A�'izK3\:W�o�B=��� 7��	['��gpH	��q�6s��g��h�����8^�M�տa�<�	�O�o�=L�d���Y3�c��ҹY�K�)%{ƭo��oփc����������u�kc��׎�U���k��œ��i����5�m�N8}��ɻk�x���uE�:�4/'\.�.�ӏ8b�_M�Ԅk��PWp�q�Gy��#������~�Fb4Ѣ������vh�����OW	x��� ���	���C�CN
scQ-�:����F��_�4}?�v꽨������Q��(�]������ܬ��a�	w�n���}N=1���p%2m�sJ�P�������<���Qf �r�){��b�t?$6�k[������n�f3����_]Lw�x���ܜN7M� /d������������d�1'�^GW���m8W�:�]� T���\\iN����:-��!�mb#������[���iU]�i�~1�Ӧ}��M0;��27�c���>�lr�LNH{Zz%�p�?Vvof �(���f�n�l��i����P�+A(�h��>륁���庩-:p�'>o�K�]9�7tђ�׶L���+;��c,S����k�?{o+ݒ��������MR$�%�	Y!�	�,�%�^x�dA�!X��0Lx�mHz�6�z!��nJ6A����n����������Ȍs�yN�����g��Q��:C��ŗ����=��{)�v]����;��+�C��X��  ��T�[a�Y��!~P�����[P�����Dfn��˧�<�Mlg4l��.��5.�90�M�颦�Zn͛�?㯚���,�is��0��u�*�����S�"+�x:����K�:U���w+1&�ê�*������@Ś������,�f�{*�*�9\ӪKS�6�ֺ#���~�o��*�+苔t��CGG)ˍ�I�6
U�􇨋ܨ4�T��!�YO���z���,�(,��F�w�8<@��é���6����Ꝧ����l�Mқ��Օe�^�z�~���[W�\9��k����������e�t!��2jl{�̱d��jq��gx07{��w.M{m�Oرa���~��ǳ&��Y��$�i���U���v��}���f��k+-1��*�r��I���w`�M~s��L�>�/ϗ&��O�m�>�L�qisD!6���U� v�>{hHC+���9��s�u�^��VxOA�֡]���l}�@��R������,9�,�HO�z�� �+��^[xe�����R�dҒ$܍��陇���˗�F6]�'�9j���s�^�a_Ga�q-�_�#ʫ�"fD��@r�?�2�g}�O�t�3T@��t�����0��^���$���;O��~F��S$���4�̶�5��u�N�(��t�������"��ێ����N>7�&���
���Qդ�c�`���<�2΅�̱�a�t>�����Qp�Lp1^L[���7M/g+��.���ΒpC����G��r$���&ċߦ�%ұ$�l�T�3�m�f
�l��֝?��,LY)��y�VUW��K����8P$�`�K���m�=oΪ���I+9Rt���פx�
]5p\�O��a
�jW�$GY�M�E7��;0�=p�������s�{�!��{�B�<0<�y��2@{������1�q��8����v��c��+n�'�m;�{��l�)�zBJ�$1]���냶l�~䵯}��G��wo|��ޛt��$k����x����B+/��IpA�0���o&�u�!xa��x)���̏C��E܏Dtw�����"Ff�ÀC6�n� o|M�w��\��Mw�@��������`��g��)�"�9��1;��>X���i�Sz�շeg6O��{ ;����s�p.Ϲwl���' re����!�g���q@kl��i���c^T��}J�7^\�@_b�����x���Ɵ�/9���>1����j�P��w̷�@ڦ��ɔI��x닟$ܻ��^G����"y�(�
=I��'>p�D#�vG���8k]�,؝�d�3tG��X���,
�Shâ�������X��K�ϡ�3�6m~��%A��ܖ:����=�jAL:���pش��t�S�ٝ�9�襛+��b��`���Y<��w�oO��	S�Wg��)d)"-�w�3�9!g��
;��{�<C�4��/���B���=��欒O'iM[Y�}�s�WaET5S��`�5�n�P��]U�i�]�{��/i�o�q3,�O���m5����Fg `W����ʼ<ۑr����<���������Ǵ�=��>�-h�}-�-��?/�n� ��'��]�@�0\�KU7��L� A�{ߖ=�����y4Nl=�hAˍ�90Ȍ���g�z`�դ�Z�x�.�\��}��r�����N.��>�a,�]ӛ�7�3��"�lg"��;<o6q�������^��D��zQ�e�������ߑ��n���כ���A��*\oę�d�[�	 ʠ����#�V���!bq`��v�m��\E�	��*�;�_���1�i#��(8؍Y�=k��q����Z�T��/N��DU���yO��a�>ku�X�@�-�ecJ�u3e����_�����b˫e�-�
vX_hۍ�X ��B��A�N�P�鳶N�lê��7��@|�������붬y��<�%�-�tm�y���'ܼ�6ni�};2C��G!6���.���w}���[�Z�-��M`�g\*�堸w_���
R꧋�%�6���X�M�oD0�ղ���p�?vvG�����>�<f$�@�CKc��������C��
�#M��#��1(��]bF�|�uG��{^Y��E��H����\y����B���:���.1}���t<���g8{�k��a�Mb���Uxyk.�7g�%
[�X�X�v6�*|���<��ꁹ�S{��\�l>��S�D0��^�1�[1��2v��y*�c-�����>b�z|����k��R�\3
���u2����*��RrEY�����f���I Q%	�mS��% �e��َ��ѧ��c�9�8,�y��S�F��3�ځ^B��n�Al�s#�{Y�ٸ=��O��`A2�'��Ad5�Z��Ս��������MT�x3+�4��ؽO�`�{<V��+��{��~�Tg^�6�YY�m����g�fk�S"3��x1����(��A[���J[��fhg��	��Q;0��'���fz��X*�KeI�з�k����%��kA.N��5 �y�ʝ{U����dچ��x��E��1ǎs�ċ����ǌr�ʂ�\Z��<��L|i���-h";�zə��N?�+�\�gtj��J٧=�(���-ء_ �re�m_���O�2t�Y��m�<���n�����5{�M�Y,�]����8���(NI���Y��r�Vp���74��h}N-�h(�]�נ�/d�Y?���w�����*s�$ˊ�~����г���c�d&ѧ�9+���6�Ud��2��[�sl;-^� u(o1o#m�!Px�Z�O�������9&fA�aK�z�)僅X\��:�HCN(�Ec[^������WV�4L�N�1�@�Yf���`�m�	�X���Gt,Z";6/N��d*��c�{e.YJ���>!��&u_�giGW�M�iv1�,c�",
�D�&=�Oڦώ��q��1�'	��eӝ^�"��¤��qAr��)��R|��/&����a�t�!_t���<y������x�x�
������\'�8r,��2�@�>o�!k��Ђ�@�Y���:}�8k�ǲ�t�^�8l>�`����%`��lh���:I���©,�#�)��k.�����)Y�a��[q'9�c��f�9�7�N$ Gm�}��Ǹ���]��Ux-�ua���SIɍ*2�7�� t&\谝���C����N�L���Ɓ�<��c	�m^��9��|�ry�B�8?4星���eI^���d��[a��?�>Z7ٴs�Mzgi�a!b7ca��HC��c[�K�G���3�l{Y���s �^ż���Z�y���L���7I?%)� �L:�{���X���U^�jy8ǺMK��	�ù�w���~���q�����)�A��E1X��wǩ�t0���s�3����؞ePx/��^�@�.vڮeL�ڼ�{��{��>�0������N��:V�v��j��	�����C�QՇ�Z"X�}���	WUt	=�N����d���c��\��:в�	,o�W?��7g��#;�������Z�{�(�V�y�#d����L>��Ա��g��S^�_�V�A�'=���zϙ�~�p��߶aP4��Wk��[�Y�߯���6�g��Z��o�C����-�i�ut�ƺ�r*�՚ʊ�]y6����,b���n'V:�~�������$JN��fA�o��xw\��[��i�7��j������E\�0�.U�w��}n`�	����K�����J�2Y�4�Q�Z��zlU���;�#h*���fw���Щ1K:�)"���z(o���`\F�CUL���{�rL��䷞y�3
���ط
N��⦵�Ǻ�q�	K�y=;�l�m���я��C�Ֆ�0�[OEhW�
�nU����J���˄�G�Ru�n��?@�1m-+��
�a\7��.����
�p�d�zA_�ߦm���YQ\�"�x`�ZG�;��kjB~ۢ����Y�YS�@���uh����w��7b�d\*����e�����]�P�߲��ꌺ=�������A;�tX؈��;� Tut�`�n�@Z��-�EdVU=I��CH�2~�-@ېc�K巿-��f
J�2i|?�l�޷y�g�:A�`���-α,׺��,~���,��@h��صƥ�pP�#��\Y���w��a?��+��?�g����/��Ne�Vh��<aٺ��䶜v}�S�͖sH{Ы׫�L��N?�"��4k`�2l��F��u�u���^��p��ߏ�X;Q�'	+ҿ�;��@f0JH��8pD�#�|�������=���Ҵ��Ȗ�@��l焆����3��6}O�~
(̕�Y��V�Uj����\��G��u��l|���
 ۶޻X{}��x}�L[�s��6a�,s�c�<k�����M|WfJ���t���$��U����h?k(�eV��F��X��E�O�;��>��W�r�S���0�<�s,H|��=��n�E���d����2-b�=���h�l���DK�{�,ub/�\^5N��)y9%n�����5ϸ9��x�w�u�s���5_����Ӽk�S�� �?Y��e��-�9��=����żw�]��1r�ߩ�p)OHzr}17^���Y�\�`��Y�����(���T'4�ry�V���ď���0٭����
4$Ke�$�5��*H�z������'}��*�X:��؃N5�J?
Y\��������]�L��w������4����<��\�X����%&h��X��`��9!�Y�m[�~�^�ru���L�Τl�{@�$���{�z���w�07Frm}� Ҷ�5/MO(ڸ��� ���z�����gP[v�Ԕ�[h�&Ȧ��beU�]�l�#����*�#*I�3���]s�u˲b秓��O�K;b�y2w���q�ob���m5�c�c	+�����6�0@;h<sP�S�}o!�zj<^���A�ݛ�7ֵ����;ƽ�7�� �����bL�?��l�(��Z�8k��E��0�9������֏'x=��G>0^[7�8E�{q/ݷ�ZA0���Ƣ̓��8���G.ņ���݇�/�/lpR�lQ�u�wl�.���i�x�p�/�b�/�I�r0W�0i��e��:��dqSt"Qy.���.c%�7Ϩ#+�GM��J�_�%�S��4����8����7��8< �z/,=g���N��^]zm�e��o��G+�\^p��~��y�����5_s�/.˨m<��O�s�l��BϪ��z�w���2��Vhq�H!��t�V �}F!�	$�z���$�^ ?��у�#	�R�ه�Q{٭+��Tpᵂ>ɼ6d���� �&��O� >�PM�T2�t�'k����(U�T:u��.��Spȕ��X�g���lC瘱eCs�.W�97����.|z��8�y6��9�j����5~�aW� |�Ƈ�>��ρlN`�ZF�S��ߧlN�1h}ˌ@���/;kA��z���#!�mQ[!�K%�c
�a�i��/U��c^�x�uE�H�]4ɦ��<t���u,�q�y�T��Z��"u׎���.I�x��.b��lEA?�	����D�s�6�h�m;U�h/~qv.�]]_���}_VÚ \���P'聐�@����z�2MC�я��٨������tu�u�^1m��`7�ش�F�;W�� ����5��#�j���(��Ƽ��&���4t����K*p4=7T)$��i�
Gac�T�ź�m���b%��9^(օl/^m��A�؞8>����ۯ0�wv�Q��H��a��FӸ�u+�u�(iP��:�qZ�oT�)O�GH��B������S�"Y�da������5���%֜4����F�Exm�o4��ru�gx���4���U�#]�0(���J~2Ƴz��E�X��EpB�![�����̦m���=/O��Y�i��U5xl,<&jY
���ό <���Z;hY���2H�vS�z��\<��x��=����h��4>�Ҳ⳶<6M�$Q=e��~_b���Mߋ���<;{o<x}̦������ �~�0�#
�6-����{�ĥ���_�~mG%��]?i�g���2�G�̟�������J��0���ec��_�H���j�!n�h� Q�qw`\i"z��;O��RX��#�
p��3^<6NR��i�ũ+�(o0`m9��p,@�{x� �r=���;�'�^m�����E ���#�qj�ٚ!��ٲ�mP���<�|�6�k���>k��={�u.�q�㍛%!1�c�#�?-��_�_1����&�E|k��� �5���9��]�+�4�S�O�**����=~��7��7�Q|��K�A*�u�1�t꓆�B�ځ�� ���Z�^����y��ݐ>�v�@��9ɲ�\��ݲ0�+���?�W�[����Ff�u�Tfo`�
~���uxF.�f\��=������gh6W/V��}�,�k�j)�	r����b>{J��Te�:���Gd��V�1g�ت�0^�|��O�B���\:^�&����ʦ�/���2�yO7�>5�;�K�(ՊF ��xNai�Mus��� �2n��q�@Ǉb� �̘���*��k�mZ��k~&����A�cJ�qza	䵜sSO륒����ʀ�x�vM���`C]L��s`g��bO�!���.���f�I�4�]<�0����E�8̓��Ƈ�ϖӱ��:��<k�{Zl����Qٺ�eH9���I˨1 Q��p�O�*塮�s���$��{��v�w'�.��!��*]R�q���b�S�4 I�36J7�q�*C;H�E�ֆ�L�H+�E9�䎳*�[۶i�W�:��뻚��u�9��`��g��B���[��G;ح@�@�X/�9��n��s f˥qX+�\�2c>0�>޲F;k���ʡ�-q��«��-c�-�̶N<�u�3���{�~��V�z�a9��ټ��?��z1���G��Wը>�h��9ү*'���,���]��v0��BI:���Ρ��C����}e�b��V�腏�)��X^��ŽX�K@z
0������q�x�qm>Oɛ]�+�ô�z ���կ��v�S��?=^����m����u����Z� k�ꁧ}�K�
�W0�H:��s.?^���$'��-���u��ې�SP-�N�r��?�D�kx�|u��K\����j��	�����R%��d0&̪�>Ix=v��󦏧b�ۏ�m�+�����h��tl���a���mt��z643�v�A�I|���Z6kY.N/u��ν��� �+ �pB�}�/��A�<��:�cI�b@F>L���5h;�au�a��'�l�h��a��n�f����&�v-A��p������ڶ.0��X��qx*�kO�	M��H˜���n�ޝ��*�����J#�8��|��S�A�u��k�nF��
�{�Jw��[R>->TL��WD���g?����xu����u%6�U�x˫��Zv�uw"��pCE��^��k�Pu%������m(���l�<�CQӄ�{��W)�9Ƨ@��Y��:�Q'��К����e�xBH2I8��Z�*;���n��G��W]c�F%i���+b�O�G���⾍Aا�-��[7�+��im#�x ���^M=e�M�_�C\pB��q�j���X?軧�8}���C#�wr�*��"
	���wg
-X�u}�S��6����y�|zl��}�o���xp�h��@�Š�H�A��i�4���g'F�{�3��~8q��G�M��ִ
�����#:/�jxWF3c����^�:h��8U<l������i�ƾ�ҪX�{@���!Z�M�׬��x��::�~PǾ�ڊ��:��ۆ{}��$�2HӘ��6� h��ө��Ԗ�iJ�,��T��Q`<�0Y
�D���b}賞�B�yd�(�4�;�-��%ǌm=y��Ň >WwplXA�[�������|o<N�7P�c�s垻n��
�۰���s��umM^�#��z=5�O�`�m�� �jĤj�~���5�d��ɫN�&�Dw#�9�qP��Q�w�G�2����.4��a.u�3��n?�4IW��;R��FU&��E�Ye7^綍o������-�>��z`��AӰ`d������۝���9�ȁg.��K�c�s�eN xi[ ����	[v�񺵎�ub	��Z U�º���L	�ԏ��{yY`���;���z5���E�VL�w�J=V>�-)��ѿq�2$³��8�u _��V�-�{?#��Y�T+��B��vȱS��`%ɠ)��7�띻�4��i.}��9a2���B�Rд=}��-�u�e�`�2|��S����s����*��\1�S�W�?�Q�B��Ӳ3�9Ae���ðc�9�j��kl[�n˕c)-���&][v�ƢHG��:N�[��u�)�A��c�?V9o��U-st���J����������o:^��\>s����s�>n֒(
>�&�ƽ���ߞ�95 P��눹A遽g��aN��w�G��{����@L�z��K���	=[�SAÂ�W��@�XYN��g�qXf��zu?�g�/a~�8��g��R���l�#=6�V�c�sq*��<�tl����$f��I�e�)0���xfu" �b�j�Ծ��V0Iw撞��Og]TL����6�^A_Ҋb �!� ��tH"=;	��da�K�w�l����6؊=e:�LzͲ�ۄ���p����r(�k<���	�1c\6oKe��g�}/OsL�~�˗�� �_O@ ��.D}�:�Ck�i�=WƜ ���
�S�i)�{�0@�a�m����'�5};�5A�9˾�aP_g�|�0��+%���A�33�Q]t����;�}��'�N�X�>����J����ZQ�nL�6"Z��������(h�l��~+D���?�zk��멤���ŖC��a����p��l�aY@��Z"͇�Hk��x�~�,c��������uF�7���) �qyB�c��/���q����\^�^�`�{9��%}�)��%��D�r�`�ύ� ��nN������M-�Č�����W$���SG�&ڈe�_\ȴQ�iN*,ڪC�SH�m�k���"yl�T��uH�%��}����J�K���Jn}~N�Oʒ_/��o������cU{A�G��%����t�;�!�u\|MPU�r@�عw�z��'���Տ�0�ix�]�����}���>��ZOsȆ(�@3}ΚQv&�H��m��
`��|Y�0d�^>�4N�������[�Et��mƭ�D��%�����2`N���&(d+8#W�}9ݧ��;��}��~�+���:��.t��I7'~z`�''�4�
9W�y���X;�SmP;R���M?<un�.$W�p�ϰ�U!'΋����������V��-p�B��g��4I�����Έ;M�F%o�x�	x��x��k�Um���^�`w�⢙�g}.�@�gN�O�f���`�w�ʅ�<���e���k�mP`b[[�w��Ml�~��ھdՀ��͛)h�{;�o�5�[���)��mf��ٶв��G�#���Ka����������
�M��al�t�u�T%�)o�f<Lʌ+�T/�Ux-g�b��+q/�����A&��-v���&�T��{I��3/A���A��n��vl�+��N�=��-�9�K�m���lZX�\^l<�|b9a�����i�xl�sBO�[K��S���ƘO?�cba�����͆1ݹ=^a�츰����l>�9�����I{�w���`JϚ�r a�շ����0�j �,:=�3㑝���5��p��;9З��������ɮ]$c;L�4Dvnl�S���H�>2>�KThe��� ��4s�ၶeT,@*cZ��K�<,����ҵ�d�}���s�vfÌ'����{f�����`���N�<mbEq�k�I�&�Ⱦ��$����:W��[A����I�W�k�T^ޗ�����B�%>Kd�m�y�x:�H:������Y�H�t`mH�k+w^�B��*]	��B��y
�����UcOI��lG�����|��c���X>/�S�jU"��`��[b�sy�����9O`͵�m�W�I��1}?^s�f	(�Nr��ϱ[fdm�V�i��׶�5�����ͳ��<b^�|j�]��G5,�7�#w܄*d����L҇�
�F3��S���9h�-P9P��;�_�
�g������Y9�b5�S��~���S�a�!Tv)̋	^Ƕ�-���l��h�m.��[ \��.9��Յ^�cG��!'�c.��)u9'Pm<9Pײz e���,��_�� ?'4����;�}z`�������qf�:>��������8T���֝ry-�Wߺ^ɺ!#KTբ�hY�,���X�O1���I^-�["��I/�1R;9�6��4h�n`iz8t�҅%��"���8����$�Wc��I:s��3�}�1�S�H/1Q��?�c�1J���S��[��ǜs���K$�f��)�ׯ�y�D����3v1�C��T,�~��i�O��>מv,��}���g��s���O�Ӷ�0l$�,��h
n��(��;�Q�e�����p�������������[�s(5���T���ꢓ"����K�Ϩ�-ν��/J�b�$jj���7���X�|߳6Ɂ
@/ݜ4�1y���p8�L���?U�ظ���ϕ5���	.pگl|�ٹ�Yfy�{���O�`l�C}[�q�2���9������-�yS�x������L�����~���B8�)����y }/�1�B�}_��!��sr�Hj�c�$�0��N���ۄ{���tz��ޗƫGO�h��
S����26,w1�Z�b�ƅ;D9ۡ=�������c��u����9XbV9F��s.s`d߱q��`��޹<�5;��3�^K�c��g�3/=Sf+�l^u��v�ش<�)���90��!Gl��43���>֗7;���'�s�C����Z�2�$dÿv2k�1��N�~ŧy����p�'g�X�gTt��Wtj��������;ow�
c��?�]���
qsM�~G�5��x�����=��exu$�u:���S?:Y�o�u�߳������9m��� h�ۍNv����aV�;@�`��cǶ�T�e�������[@�嫉���&@�A��-{+�i�����*h^_��m��`;!{G;t�bG]=|��$A��i�z�5���O�Vd~b/<���NtƨJ;V�XK�c��ӹ�C��{>=.���k�Ȼ�� ���L��N�#Vէ@�eFRbm�=�kG��x��T������cѬb���n^��VO$�����>������U�(>��j�/y�~�h�Ů���z�yh�ߪ3bs���
��3�&`�EH�@]�{~��R��nFe}.��J������5��"���<����^�]����|��p?Lw�K0�[>�p�S�:6wV^9g������,�=C���k�AS@�����=��� c��c�^�:�r�z�����qj\Gm����K,~.߃P3���d��䘞<�l}�ظp&�J��-��e����hof����Z�?��&��z��������!�{���3G
��z.mt����2��������AG�-
׊>�"��S	���-;>Nx�?��b�E;�"��E�N��(V�tV����-S��J>mQ�o��8����+�Y6����ڋ����5W�9 �`�v2��{�c���~�Ҟ�Gn&�	{��f�����c��{�{��t=��	7/��r��o���
 ,�%9��t��=з�۾�+ U�̍	����{�a�B��˵;�a]��Ù��C���*��o�\%o��Q� �j$�C���A�Ә�=s�%��;�s��R�Њ ��"��PwG�ݪ� �[�{��!6�6J34���jYb�9�ˁ�����D�c�8�:N���/1i}��r�c�9��1�`a=�����P%���q�nr}b����ܻϵ�q��syDЙ#��[��wj��������An���ʋ�U����|ߍ..��X8��x�u�7��S�mh]O�����v�H��q��'����6z̤Ԉ�������P�ŴK��^qڳ����]��a�_���jM7�k�;�@�O����]��c��� ��C�(���@�c(K����~�G+�Z�g��%p���X���씭�K�����랰�1޹�́��ցzdrG� �r^��˯�ۻ����{.]���3��V�1e��,�������2^�x��������2�n���uG,;��5U��ꚁ�ĳ�!z��욡��Ы8H�kX����m�w�G�q��H�i�����~��j��I4��"�ZG�D=/��j�޴�p*�򞵝r-k?%~�e���)��{�gb����I`^��9�k��?��߂�U/OKL��Pt����h=c����b���a^q���g9����͆m��{��9 ��Y�}���7�#�~]IF?��_�*����U�ڎs�PG���������B�4E�\�����}�����i�a�ӊyR��p��->�U[J'MP��5^�����ބ�؋F,{�G�<�x�-YH�7��bw�M��2h}�-�Nhs�k˺=	�v���a��-���m����z�סs�6����|������T�%�n���g�ۋ_�t�rw�9�5F��G��������xB�A�|/_��%%��>��+5N�����Dx)�cQ����`�a.�&�� �1�8F�b��rY{����>*�u�cY
��O����Us��O^�?}��ő���^��%v�]\�Uk����D�VsC5;�n�����KW����7���N_s�s�rZP;e�c~�Иc�K�s�Ԗ�,� ��[=�7e�6v\;(�g+s�S���K.��s2�!�>�q�)o�����T�|a�6Ҳ!`��cXG6�\ܞ0��ܻ޽9���5�.q̨0���c�G&���9K��ߌb�v��Glߨ�g�򊢗�vHex�q��*e&����J���~Ĩ���>
0���>�	���o>:��vM�C���wB����l�?�Α�o�qQ��"��J�O�Ur.����nwR��9�^D�u҈�QT������K�i^J���+�����h+����H;;+��1ay0u�Ñ5�3�s�;%��u��Zż!c��m4��?ޞ�>ur���:W�ի������L�C������Xjt�zIS�����L,'`1/��-�Ƙ߹���B�vខK��в�P�+�8�6�{}"X���p�
�g�˚��T|�?�z���(��:�c)W+����wr�ƪ�y�:0g�>.�2i���`�2|Q=��ج�=Uf���<q~��1Y,�+:yf��s>x��9b��p���k��[ƧA"���`�Uҏ��hK�m� �����籓���Ք)X��]��m��.1v��1���@%��G��z��6����c��������Iy����Q\mG����A`�	�<�ůq������#�{ݦ���,ڶ��LgƎ�ǹ>-M��2/��ܬ�˿�v#�#���ҼBS���z+��69V4n�t�D���	�}<��O�_����+@o��1=N�Y�g�&	�l��XQ7&OL���e�v@f�m�н�ޅ��1�H�ä�ي�[�r���>�(������-���9>C�A�UMf��O����zÁ2�3��M.����w�`�Hn� N��a��	�>�+��"�����"��9��yʁ>~l��ߜжB.G�rcD�a��þ��Nޣ�][L�dž,��3��L?��ZIg�0����]jƻjRw��-��½���/�W��j���7[��Ͳ��Q�r!t���^|�$[�&����`��m�ڑm����A�����K����\��e] �=+XrueC�^�yzBQ��]�x��KB}�%m�k����� ��30��N��Cz�\�y�����������S�vw<����\�^;&Oz}(wKGe�B@g(�yUE�ʰOI�B���f3Yl��p�L��2�)SŴ�b�*,X-�8��P��a�32�a�qЎ���d��gn���3���r��j��s��u��1����,`�:�}��%���� ��u����	S���a�Â�X�	k4����g��k�� `�@+'H컹��q�x�@r��/�B۟&޸���kc�	O�3���>�c�v��>��-���qA�Hx���O]bޅ�鳿�$T؉g ^Ѝ�z�C�.��Dd���=�>��������٧N�3iĉ��ӧYI,�R�́?l�Ϧl�J�C�Y�ߴtss�~�g<�TS������@[P��s�	Ox�����Rx>(���k^~l�y��:<d o;���{e���$Kg4��?���=����Wv�aZ���'�x�4,GA�>�4�^�Ј����թ�M�!p��u��T�^O��W�dۧC�}GhQ��k��\�AW�= ��k���M:S�½�>�ٖ��ڄ_\Q7�錈�"��xV ~�����[�wE\�f�ޱ��,N��i�À7�j���c��Nө5x�i���w vV`7��8N�S��-�e��x�YoP��9���2ǜ0�-����	�\����h�娾�)hx;���m��<7p&�	I�/2D�؋B;&��k����ٖ�ˏ}&���X�zD?70���Du�n�d��>6�Ʋ�ۅ���I�g5<c��ĩ՘�1��Z���̿>�?�4�6���1d�0��1P���4����2���B^�
�tvi��*��-���/Lo���o�$�z��2�ۆ\��t����O��)�p{,|.�~iX�R�"���2W^}�{>�N.�z�2kk������x�8�nS���m�9By���[G�r��Ђ��|f���c�濪���|��A���.F���?�T`#��e�0_t�P	�ޚ������갦�y��Gı%g�$s襵�ۄ{�m�7��8�[=��{;�B�W�u\�-/�����8U'7��o�a�5݁6]K��|ssE����P-O��sESс}��ױb�s��M:٦,��R�ۄ�_a��c>�Y�6��9{���S����Ѵ���62};�ԆF�v�9��A,�N9�I�[������KмZ7�_Ϳgz���M-,�"H��m���ײ }�Ĺ�{�W:�?]ͱ՜9�P�T7Xwǜ��xm�cߓ'
J��.|�����.�k�~*,p�?z/�����~g�vk�{/��A�,d��T��g�����kt( �9#�����1_�.��.��?^#������a`��;�u]��d��v����"�'?�Voeog�O�k�2`�9����=	���p�aHj%k]æ鏩X}�{A�P��*��nO�>�~���
��N_?����8�T��"aT<��=�����:U�硫��?1~ˌ0x�~{����F=v�9&�՟W���T��>����rSQ
��?��}_�lw�z��k��ɏ�^>�v��"W��l>��g�G��Ə�;7��	��}w�g��l�?�k����������N>c���67f�ޒ������O��R$��x��X���^L9�I'�*d��~N�~�p����j���v�3��Pu�|�Y[a;�TB�K�h�3#���
���蘑00�Ζ&�@�ɃǢ�]۠KB�������,w��2`�`������zk,�X�:���d�;��%v�`�#s o��)�h��w��{���
Q۟���u�q�B �kVgo��� �{V����D��"v��|ކ�{�$3�T)Z<�I\��S�u����~yp���Y�%�_�VګTD�"�p����[%�4�s���{}��Y�sjy���헭�(aA
O8Mw�J���+�g����8����cZx�}��������A��'Ngm8`��f[^��6`YO����i�~PH!�ú�XhlN	4l�6Km����S��'�<�g1���T��#5�B+�[�M7����v�j3k]�����S�1���j68z2p�S2�y���X̗YO��	I�i�-���L6K�~�tLb�ۢ�>�a��ϧt�KZv�Į�����;�Y���.�)6Aʞ�m�9}b��ei�=[`W�Ը�U��2���o)�c�|�oCnP�2bԧ���xv�[$��LO߷��Ə�V�qǡ�g_�z��9,S��W���+�Zn���˳���3��d�� ��\�, zy���\{��{_ﵝ�6���7L��9����M�Yꢦ&��b.������|m%�<�3��t�=����B�^L�떢�`/�^�g�	��r|H�NC�[%�1!ƻ�S��ъ�����ƃ�H��S!T�p�YC�@Q�N���?ip�Y8�t6x�Ǔ�8Ne��Bb��b�����i��&�PzSo��g�l��^G�Ma�����>�3���iA���|���x&57����o�<��^�9p�z�Wn�!>�-�r�-��4�o+0�?b}*)����1kӕzK��We��`]q"T���G#��c�*��w]\ی4�Ԁ_�ՍL1�q~��Z\+�#!�{��j4�p
��*_���|jU�C��6w�xZ=3ɳ���2�M�e����1o�	-��� �qJ}���4����>��ɝ�c�V�`;�^<�;Q(p�u���x��S1����`���qy �=�N�}zB���1n��L�.�/�3н���ZT/��9P�����������v�&)�Hy.V)�2�������o�y⋇���BL�cGk���ݏ�I�@�+D7/��uu)>����5���+����Wɛ�I�ρ;������]�%��b����wЖȅڿV�}2��OT���~��\�j�|����w�c�r�r `�m�v��:G UsH�jJ��±��
8;����
��LC��OA_��|a�y��n��.�m�y�սZ����
�'�6��ۺ��yV�˜���v�s�P`>-�{B���lyu\[#��|{�����=�L���F�i�}"b�y�G��.y�7'y�������ٌ�,����
���� ��}�ͳ8�B%ռ���b�OԱ,( +��xf�Y]ѵ���ܑ��9m~��-`�ŃS���Ƞ_���'7eU���04Z�Ȕl��FW��j',��A���dV_��t��hzȖe��|Ep��m� <ꪞ��4�=h��3&ͫn���i�h@̋�K�z��c�@�%z�n��j�Fˎ��:�GCj�v�.m�����?Z�h��q��A�A��Ə�Xs�C�k��<Wܴd�$�KI��!�@>#��qW�����6
�����v����*�c��[�Wrއ�c��xx+�Z���HE.���\��[�U�ۊQ;��-Z���hs�V>OO�X+7��r��2��i�@>�pzF�2]���Q%lP�l���$��7�X�<l��,����Yԛ�ؖ��%&����������j1��v�RkiЫWB;�m>�w�7��ʵL� �z��aa�rX���x��2͹��v� �CN���k"�E���{u����÷ܸ�{�
)���ÚQ�C���HP�/�X�kQ*\p6ҋk�1"̙��E:H��:��_�Ӷ"4����,�r��q����;֥G{����D����ӌ+ڀ�#w����8EJ��]�
��>ͧ�gO�����h����`�"v�S:<��LY��9&j���)ū����~�i���cw��Og:6��`�|�2c���� ��v<ʿ�O0ݜ*
�kg�<���L����G�ƂƏ��
C+���G�l�s��W�Z+g�=�ǝ�\���1u�P��E]`��֥����:OV=��P��!��P7Y��V�hp��{�V�@(�`��3`WU��w�!�*��S�{���ЇC,����A�ϟl��x�Y�H����4i�Z��`��㠲�q.X�{�cy:0<0�@�.op�,9<�i��?���U�t�i�M��}X�bi��%�cAٳ$�*�#p�E8��o�{�����s3��4�^N����p[�d�Q�z�����8<!��G�*��" p͋�MKE�!���~\kTU��k?�N�*!hc���A˹O��S��zM..d�[��Ӊ���T+꼢ݪߩm��s��Ȳ7���4*/L��W?�zΥpʳ�̜��c�K����_/ش4h���ԉz��	1��{*��?���S@�c����;Ǿ5}�y{V�L~��՜е$�#
2���>2q+���7��G��E��x��O��˻�	��K���S���uG<͖5	E��?OU���ۂ�������|%�3�ӫ��cM�B.�O�F�h�-�vӸ�Y�҃��}��[+�|���Kx-&���  ��&̒"�������;�,}y�s����m:�ɇg��V]��R�x@�u|��g�g=v���G�+�]�;v/�?{͖ˋA�+2M9��5���aܞN�;�D���ű4��rx��w����E[oC|N��;�o�ۜ���9���re��{�{(Pr����UΛ���f|�^�uLǪ��B�[��Gߗ��Z>�M�kxHK�u�`�%���btl����^�ke�B�<3�}Za�iO��N�|I�Fs3��gl�1���nD@�bx��]��l��A�esj��X�E� ���� �şˣ�n���O{'fYƨB���5�_wf�����b{�qX ��6�V�̥��dˌ��i��z��{fNh-�|���(���F1��x��ɩ�4���WW� ǲ*�w@\Z>�=mz�_wϊ/�L���2�YR%���"�=tR;����v�,V����3��T��[�ټRWr���I�'���8�S�f�a&l4��`���bsr��L+)V�<m?�b�(L4�1ݪM�<��9Fvʠ�&��
��y�g 6ݹ<-|;$�p0��]����7�m��Q��Y�9�W����Y!���ͱn�.ZOh�ZVǂ ���9ǈ�w��~��qzVj^�z����w���gi�c�����#�o�[�ao��$�=�]X�S��ر0��*�_O��8)#
�=V�����&�S�5�JL�������;���z��7^���鹧}}MM���YE{|�堁}W�!T��������ϭ�=�=�x��%�ip�O�!�Z*��]Ke6U<+�����e���A`��uKu�V�sz�{C�&J.k��`���k=z �҂��ݓc�*H,��� ,G�oyTv��7ډ��is�Nӹ.UH�)�2=�K~��;u1���=�O& Bi����3�e�x��9���,ZF\�@�E��.��:��RR#��������Q�i��*p�m����gkˏϪ�ͭ� �W��tP�m�uLX�v[gض�߾m{L(t�7�3�����QQ��[ ��p�u����4���3j.����d�;����P��Ѷ{A��k�.�PK�V�V7�����6��z�,��<���*��E��i]r|�Ѿ�2m�'���5���SzP�.�k�މz^u�U<uϺ�N�-�,f��d�;y�o&�q��G;5��#� S+�g=L.�jH;��=�(~ǿK3 L+w�^�;�����/ǔ퀔O��[��I[os�^�BӖM�����2d[^�\~rm�e��G�ˤ;�9Ӯ��!��}��9�j���������L�K+���Y��Oml��O��}C�Q �_;=��0�z�������8m�{���I��d+��\�+�;��wZi}x�$ӥáO��p�I�Z��S%���w�s�b"5�9q��&��O&bѦ�}��o�j��^�(4�����	p��b��eT<���ݛ��;K�m��.{�j���^�a��t�གྷ �iX5ENڿ����y��;0��[�g�n��S�������8���b~�Y�/���l�)Δ�#Bs,�N6��;�o��޳6�4a�E�λ����^f�}���YSW�I��v�e�J��r'�|d����o� ���ʧ�~Qv�l����X����+��fԻ]�J��Q�U�9�I�v����Q�/v��N�(�0���]��a\���i#%5�w�Xl�=����w��\��p
�c|v
l�Ҡ�]?��F,͏��)�\y={t�c�?L�	a�@��|y�̧�&�M��N�?�WL���㳹��\l>lp.	M����l���;�����	��r}+�{��uĐ"y/7�Ί;����� =\=��ԥ|���'�6��c_F!|���A���!��iV���jԿv�.��x�0���/��N���%/�l�Z�����V9c���i�]g���7[��/�*vƶv��e{K�М��2L/xzi�/�9����nء�c�sy� H��t,8ye;�^l{.	|�֓�fb�2�Ǧk'�|*PN@���?4R��t��l��e�>l8ӱ��g�8<�n��Z�X�<�X�sGt+a�r��V�����3��u�1�V�5�GO���<_�먲��4���h
��|�.[�wUeb�m�XH��ͳ�5����1}���i0/�T,�֫�:���۱х�r��;�Ԡ�9����2&��/`��bi�>�g¼�����ڼ��D,���S�����s�M\Y��s�����k[�����t0�k�3����뵽���'s���z����%���8�r�+W9B�B��i|�l��類���f�O|� �]-�6t�'j�Q`df\3 ��D3����`�.r��[����ʝP����iJQ�-��vG��9]�+�%^��,9���W��;q[�R��b��8��Cb�qC?�#Y]'��j5�+��4$�ƒ��M6�?���~����X��ǿ�)S���,`O_�a#(`��r��!˴��
��2c�q��8H�]�ȕݫK�����	^4_^9焜7Z�^>�Zn�^��x�n�n	���v�٫��Q�M�;��xY.C��*�Ґw1
/���c�R��3��[%��i��)�83(�4#`<c�FϾv���Kb�~�(y-�O�߭dW/�q̀�m�n�5#ѯ��-��?�'�U��{����Nؾ ��U�z�ߋ#9�@�,�ꑁ^2�΢����� �˨��{w�F�N��{C�xJ�h�o{m�yl�~�0�y�Q�[fa�;�~���wB���rf<�c���ű
�$4�B@��+cN Z�����[D,�25�g��տL��(����~�M<��D ?֤ӫ�nF�x�Q�����n�7'�z� ���~=���)J�j�q�����Y8O�!-[F��<�_�`�c`�I|w��`��������߸(��Wtv��ޮ� �o�t��y������>�D6�2<Ð�kҪ�����ćn�ʈm���{�~2����
����H�*[��?\oycĎ� �Q��@��Y �MK�nP Y�ꁡB��-.z�Ȃ+Zo�	jte=Zi<�y.FN�$�_�~W{rTm��C����k����ƥ~��}o�����N5䁛�?���f�=���{;MA��qH�l�!��K=����Cj�/�{|����
8�E�ζ�]��g఍O�x]���>��/u�mY9��Ղ8
j�cڞ���d�{�^�T��}1��(��f<3 ���r��m&����o
9�[�}�P1�K���]oiu��6_J��W`���`"����E����ݿ8(>{�^��Łd�R�������u.X�i�S�d�:�83mV����Q�a �7��s7��[�M\���;ű�T>dY̔i�`�l6T��Ig�07P�CY@B��
��F�/���B�c�9��g���}2��c�`:��x��k��{K3'[&l+oV1�e���6���;"0��!9��nh����_a���>�ǫw�~n�X��y�g��gI���w��r�Q����Z�맶�V���S[���r$u]�Ƭ��~���H:��A���z�v��������ɽ�;t����!�����t����kZ�=���ӟ��̓s*ojn��Qt��g��Q�kh�j�r#:2�
���*�$��^wN��)h �i�&�y2�h&j�\g����l�c�9���Ə!'<���7���k�97`5N̗�>r���qPyؖ�2�� ��$O&^�佼�g�t��Y�����g/������g����*�9Xa�ҧ
)/����[�`ǧ׾�}�s��%_]Er��E�����\��q�a���	��-}�◧(����͗D��|z`@��BN��v�h�>������G�Կ����-�U�w���[������t�=�����?����������:�w[��#]�N�/,y'6��o�}_8�F��a���ϱ��A��~�:���1���`�urؽ�ls�@��	�W�V�KÖ�[�,s���Ws�.�9��4�OY��&���P/4�dA�϶�)峆��SA�
V/X6~�;^�m~������i.�3*�嚙�����ڣ���czm >k�{V�̹z�2��s���ڝ5�7U��*0�=����O?�� �� �o���,��v{*���&|���q<}�u[kf��Y����_�
G�~�>����f�(s�V���Y�"qY�Ŀ��4E�vĴ<׺;�`X��),&�:r�Z�t��̗�)����	^�7�0�hb=�#�4x�Y/�Xe�-=gLL=Ad����`µ	+E��6�t,`�2���{F�_�f��'�s��։-�}��crm��B�2�2��H~4��iWi1��ƷŃf�~�r�mX�=�D�OŪX�oKO���1�+�E�,|��y�Z_0��b��j`T'�
��Ç�È�"��g�ԇ~(����c���l~Β�H�\����p���%���g����?;O���v�L:�����xmP��΀L�G��zAM�E6��Ͼ�	�����U��ʁa:�2��[/Ϟ�[��w?Wsi{���m�;:�\�ʕ�c��n���5/($m8��z��=뵯.Bk:(�?C� _�ϕ�Ɨ6x�Ď�\^�xȬ����|�����Q`�=�j&�ܼ�Y����� l���b��Y�aw,�X���.}��g���wM/_���77�*�i�mDw߱j�I"y��x�㝻�x�h��XݰU�[v� <xk���e;���Z���_��%�ֽ��Tq{@ɓ���s�c�t�X�r{�Z&`>0� ��������1;��sN����^�� z��T���fZ!��A�a�W��v@�}N�=�D-���U/���z5�rydצ����i�����Z�a<�|�������b����{�2���m?�S0ִ���~�8����?m[�j� ��exje''ju�6��xr��<�u�-mwR�~I�o�*?/ނ�>����*�]^�-�J�Xl�O�z�;�ӧDϟ?�w�5H���>�������l��'l]����vʈt��BO:sJ�JeJ[�ߑ�'�$.Sy�`m��XFnz�� ��5��z�hl�V}㥕�)�T��Z�� �6�hvv�����~J<���r����i��8lGk���q]G�d0k��-��qmYH���տjE��E�zͫ��ƁM�}���oz���&�g��v��m0hh~��1m���|'8$溬���m�꺡f��C�>�R���{H^X+ �������ܻ�o��;�|᭯�?~��������}:{����q���]���i�5�>��6TV��{$d`�M��ɪ�;wyG��Tӿ���Gq�740�'v���V{ވ�m�̡��T�yf��TT� � �Q�(G��}���㙞# 'ƞ�8b�k�-���HU;�߆�+��O�_R'���Z�NĚ��O~Ɏ�^O�{}\ǐl��nu�1��*ن��m�u:���*��J�d�|���`K9� 6O�HH���}fd�5ڀ��Va�绶���v�RW�_��edd�n���v�K�Vgaz�U �^i��u�'���ΚT0����w��`W��w�5���E���V��������`��m�uT���m'�P�L�m��>n�N���z���~�5Ɇ�����E��C�~۩!D�7��N���	TUL�UɈ�v�O"�#N��Lg�}�w˺kSEL��a�Rᄂ�J�ܥ�'�g ]w��:�F��W����
���F�q��w�R��h�]L�y@k>�C�x�H*�
}3|o�Cf��jf�:?�1�5ĝ���M����M���|�G��<�\�ω6_��2��/�������������L��"}�'~�>��Ho\��7�tW��A����׿������9}��ߦ������WE���+:ߤ�5��:H����+~��paу���|m�w5Ik�V��"t�uU�Qg}�¸�jx�,��7��Ȫ8X����2'��j��e�F�L�������3r���,������=�k��x�Z���� ��ŉ�W����6�Ӯn$�%�54'���X^�a�Z��ʫ�`޽Y���qVhˌ�E�C� �
A�'��'�u�������u��ߑC���/�npc!�E�ax�1�~<��m1Z@>X`7E3�.�*X���i�A)MT�h�_��(�|8T��09�p�Қ�,���y�b�]��UuAe����K������F�=}��~��������t��BZ�nn�½�������ӏ��3��?y����_���������ջ���տ����!n�߽*2���	�w�}N�:�*?�+��a��7�aF{�uq��55�U:+�����;0��T��I� ��7T֯d�լ_��a����p8�4\W��|�w�FƎ�l*��%M|���
r�N��BJ'8��ٻ���nb��-�Θ�qj����Ī��4�밌|BP`�E����.mc�z�����J�լ~�I�q-�
��33�����i �Ct��u�������� ������$T�������x�8�6<��eR�P�T���\6Nc�ͪH1�s�����?ROiş� ��,�Ӡ���
���.�j�bb^%Ug�,�x���W�`,F�=�v�����iOu�E���a4M���2����ϒ�agwя�1B~�����z��WJ����I�~k>mw��0p)���b�qww?�A�X��Tœ��R�ZK��?H��r�y"�j�e����Q��~70�gt^�tѲJ机݆?z@�����[�G/ߣC��!��5�Ń�p��߻�G�����?����|�_�*`�7��6�]��o^�]���Z�L$������?������}��={F_8{c�ĝl]���x�~����[�	y�����~�g%��o�6�M����R̠��U��=��g���nj��d�ބ��+j/�	�9��U��A�
�T�^��ȵ��dZ�)��}�723;k��xn1S�ؙ�w7�ɞ����ڬ��W��dxz���J�5S��W��:�����F_�j�lS],`]�{�`�����Ǥ�� փ�2���Nb�X�v=����wu�g_�"�����Q��/���f��u= ݖh�޸����q��(5}�G�+v2���~����<ps3ާ�^�x*�����1.�6To�zk2./6�?��g|�����9������s�����������飏>
�����o�{�G����J?��g���&��V;�>��ggtW��A�>{�����+?���z�y���=���uϾK���ғq[z��}j�����߄:�n��Þ��U`0q��z��|�b���'p�7gabpޏ�{>6�J�4:>���=B$�f6M����7l��k�n�d�u�1KN�B�X�q%_o!L��"����������H�I7�8Џ�1=�f����qk��^�O ����p�£'���/�u���5����4��~�|��B����N�!�Gw�<��\ kM,U��g��s�a638֫�5�����2	�ĤjR�%��qF��B��0�+#��u���L��Ц	�:�yL����	}�W�f:�ȥ�Ǥ���4�8fƩ}�L��Gb^���١�����
�X��iڞ)��:Lڤ�^Ӯ�3�Ch��R�V�g9�!Nǐ/�wm���.,�����nS~.���A�����U��_�t�Q`�j�g���{?|&^77�.� ��{���f} �������ۡ�ޡf���;燏�;��]�8��B�����џ�3?G?��0K�o�;�*�U�w����l��O������_l���ߧ�|�Ǆ��@�����w��x��3�����`۱��օ�('-^_��݉�#a)�"���>�N�kk�XmDh<��	+���V;=ϧ�5�´l�BW�����7�s䀝12��ސ�u���E��vn�7+(�i����<�撞\���f9�I��㳬�֑���O�����m5���3������ +UGrm92\�ǩ*�dxJ�ݮ�`��������st��e��5��^:��er_���4�\&\���U��e��Q̷����i�8����ıɳ]g��bߔ�m�@?�� ~{g��Z��M*n♷�����h����t}�R�c�����k������ky��������P�a��tqq!���3��Db>7e�L\������~�7����'�+��+��o���Gޜ����k�j����/���P����M�-�����w��}��}�>w�o���{�Gu�#:?|wX<S�/�h��v�.�R��[j�#g��^nC����/�PaOw���K:�#� å�qJ�K�;똚�ؚG�����ݡ��!�v1�.������d�(X鵭5;��8H������@�Sv�T��.D[u�@����<෬Z�gd�Š��y���4+p�E_|v׍�Z�W�D�G��֛䵘z��x4P�^4_ru����\��}о�qZSO+���m�� D5 �q��߂~\�<*.�Z�H��2�oX5r�T���LmYU��B�U?!����Q�`P�Ġ�Ok1�/E��:zu}!o�F��(ۛ0��h{�fϞ��i�����xC��[�^}H���f�~�BZoH������6�9uUK�ޥ�� �����=:�2=��w~�A��G��o�/���/�_��?O�}�6�,ଥ���N��7��'O����\�+��o��H������eo���O�a?���	��y����O�״9$���U#>|���Y�v��q ��3��O�<���
@Ϡ/~�V�1�Gts�~ ��X�����&���v�Ou��u�@A �}#��^}�� �i�`C6��� � ����@P͇걋z5ċ����
Z��*��F��\4�늃~��*��E��r ��<_���:�3.OТ�T�:�*��PO�L�0�گ��1-%Xo��u����{z��e0�Y�os��_މ/����0S��b���w\gѶ��b����'-���0�3V�_��כu|�b�@�دzq�^uaV��1�B�?�L�$���Wtq���9�23]�2��8^�>w~��/~�t����?[�lna��g�<���{���_��	9|��_�գw�}���ax-�O�9�ޥ�jK?����݁.���7~�1�ؾCe��%>=�f��\�a��葨w� �؜�;l�j{MU��ͣ��\_��a��yf��w�E�C��{�~y:� PY0����D���h��zֿ����EPd��	�]�����S��@kî5Xf�m�@���c��{�ط�^4�����a<�t�8����'ƅ�뢜WL��UAXV|j��@]*�R��m�'�ԓh�]�c�H(�Q�ŮV^�x��v���TUlѰ��'��>%I�XI�H��q�g�c�d�}��z'yz��"tV���^<{@��/�7�ًW��|@��A,u�޼Xs����0#��X�Ś���k��./ߦ]����kZ=n���+�~���#z���/~��y����xW_�%jYE�ޝ���;����x}s-z�G� /�i�6�����\�ov������c�y������D��W;n�`��G��+������^�\3}V�}*>7uGPĐ��{A�e��[7y�Z���s��Y�x�����w7�iD�B.���Q{�����}��y����k�*�P�3�ʷ����m��R��5�=��;J9�̲u-��7���(��M��鞛�;����>�S�������ʗ�
왨w��]]?����}<����ъ�����ҵl�݅w_жy)ۑ�|�}�K_��|xEo��foӇO�񞦟���
3��>���<����,����������t�.aZT|�6<�ߟũx����4��
zkC](����9�@&Ӯv:P��-����Z��m� �+���D���=��+�ʂ�,\B��'��߾U}����!uHs��� d~.�a�'e�k/�0�;o�M�6�M-T�o���|�>�����'�/���)8������N�8���t�E���..Y�@�܉w����=~ ����|ʪ���z�1���#q5��_>��;�KO>|B����ӟ�������g������wh��l�����[ϒ�%�� �o���H�C��?J��(�շ���d��n�b�|�!ʼ~���]������M:��Z�W�5���~��a�$�~wN�?�o-@�����·��J���9�g��Y��E�w��_�Ō'���\]����u�H|���ɳ�����ަ�o�*)�����ӟc�����s��?�:���`�usMO����W�w�K�ý��n��V~���|���<�������t����O4�&�=��ش�a��Rr�5��D����� ^ѳ}��Z	�!Z��)f�* >�R7tQ]aPс=s��t�&T�5}>����]��~�`"��C_p�����k�G��%}���O�$��m�|���<�?�����S�fM/��.^�Ak��;�㽃��~��/��?�=xDW�ߣ���=y�C��Z�;Z=Z�\�
���E��U�l���10���8r�"���F�*�i�h��n���a+��_?��}>�����������?O����[?K����֋���ע��������7��
�~�����ߕ������zl�sy�Sq��ˋ"��۱/���I�Σ�(�[��{�sV_PY�y�[�ľ�(0�:\��-�U���L�<���4�ެ���` ���5�F*��2�%50Х/�0u�
�̼^�E�5,��HT�b0Tm#��l��[�w׻_+��q��u��W��\��#�|���Y�m����8�~=7
��-g���t�d_�\É�Y�q+ꐻyj��öe��]5����� �Af�/�;��Y��F��mV�`��߫Ѕ�8��F}��~��`���i���|��  ?� ��� �B B��B} P� 
y �zH.=p�    IEND�B`�PK
     ��/Z	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     ��/Zd��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     ��/Z#���5 �5 /   images/4ae07c11-480c-44ae-b2c6-f8186e930d96.png�PNG

   IHDR  �     ��?   sRGB ���    IDATx^�i�miz�|k���xϝk����nw����q3D� ��)	�
	"���A���
;b`!E!&1v�I�NwW�T]�;�s�=��yX��[��u��J~D�K��9{X{�w}��=��>��)�;�,����;�,����?�P?��`g��v�Y`g��v�Y ;P�;�,����;�,����;P�;�,����;�,����؁�� �Y`g��v�Y`g��v؁���Y`g��v�Y`g��v����;�,����;�,�������;�,����;�,�� -��>ލ��v�Y`g��v�Y`g�(܍��v�Y`g��v�Y`g�S�;�,����;�,��������u]+�X���Җ�03����@��Ο�����à ��y~���Ls�wM�y.���N�V@����������+�*�{�|oR��ʣ=�������xq���ɺ~���g����(�jm�����{�����c5�1��R@W�.[{A?�󼪕������Q��r�1�(��~m�O���k�}n���m��}zL���}P ���/�#�ݎ{����i�>���<�����>�l��!6��ڌQ���x?Y=�{;��[|��$<k�6�n��}��x,>h�s�~�x����?0��I����Y�9$cR~]7c��8�84?�q�?n}0�Ձ��nT��v��z�6&�177�a8F���ef�uY��d򡹗{%���"�,۸VR�a��$�ͬ�Z��1Kߵ�ʷğ����L����ti�]x�e浕f���ꄽ��C%�P~s<(C)�����L�ʩ��u����U�u
@���U;UM!�gJ�������'\'I�ݼ�Ӌ��������]?H�G�޻�߼��>�I˪�(ԣ˫���i�n���(���mI��ʰ
Ti������Y�E��jA��y[�u�w�4K��f��Z���@��k/�kO)��rð�$IjSY��.r��*�®K��en�]ڶ*�MS喲�J�u����J��PU��Q5j�4�ʶ��2���Q�y^E�$O캪�a��#6M�`��j�r�<�Q��Q�.��pQW�aY�ay�Y]�J��6*�4Q���iٶ�P(뺬��6K��Q�,�Qkg�N	ۀc�u�@U�YYxU^�eU�^��'E���u��6~/V����Tu�\o�*Q�UU����6K[�em��8ϡ�+�(K��x��I���ei&WhU*U񝕪jU��6JeE�����3�u�efV&���ҴTN�W�<sU+�Rfium(�T
� �2a �  �0��+��ʍ"���UU���좶��VF�L;�,�׵Q�e��
6�ʄQD�j%?�4�}�(���*\�����M����G�[�v�e_7M�tl���RU��ywQԅQժ68���.��ʒ��B��A�2��8�"���*��kUGp��4��4T-�]Y<?�(������`�0MU-W�p<]�5����ڨ���+�Q��5ĞJ�Q���i���	M����fY`(�rL���Mϱ��s����`,�R��Q)[�(`)�3ժj�� �ʺ2,�kJ�Q[��5j3I�W���󼬮se�Nm6�����ge%�#�̰ӛr<eY�*FYe����jUێ�Tu�Lˊ}Ǐlǡ����"ϭ�(�F�n��e�J�Y*MS�(K+OG&��9kV<?e�p,��K9��8뀲�4��4L�,��-�(�FY��+3�.�\�a�J���TN�{�[j�g\�WVY�8��B���,�D��5�Qy�[���Q��a�F�Nœ3M�c����r\��+jUѓ��U�Piy�����eM��=���|o���Qr>��g;U�E6ϻ*J�3��͊�n�����P?S�RU���V�zbX�4��0kv]U��(UV��,sy`^���[���a�Y�LǬy�l�N�$��)hg�7������,��*m�>P�tb�L�(M��Q��Ur|�Fe�N���Q���ZQU*;+���[O.//�˼�\ߏfW���w^\L����v�h1���u�/��M�ȴM�J��-���*�4F	.uap�l�P����eUXUY��Ǳ˪��,�_U
�a��a��ݨ�܂2L�0�(겨k�q8�Uo�a�F��,ʺ(���\��r#+re�~�&��'��G/�����J�������$�����ؠ��7�������ܳ��L���!�cX���(`6r�XC�LzC8���l��v������-�y�8�"�c��3���N���N����PV&�5�(C��ç��8-���T�`��t��8���|���#�9׭gVU����y��9���Ǳ��e��)��w�a(�G:�Q�aݰ��u�|��Ry΅�T�몺Rʱ:<:B��Qq]��W��-˂�8�<_7�}��G�$��:�@�7�x.5xe�7���Ї�&3����ե��.
���#��#�@m���Gհ��{a�䕼�q�*�DI�`%j���:-��24Ee�&Lۮ-èKM��<�4XTp)�Fۅ�F�Rq[��`���e��u�qIGm[�A[WJ>G�����m���S˵��v3�Waȍ�{m���"���R�>���k&�uMB��c@�|],V��`��3ʐ��F1j0�DRU����{�8���Y�!Kx�#�q�����*�|��j~��Or�P�]���m�AU�u�&\�˱�y�0,�2����<�v��yۖ��܏��H�L>k&J���=������A��R����-�$ϸ°-���e�M�$�ks]W���L��eY��,����<�]׭|?�����k�
����i�2�jj�Fmf]��g�i�r-�����E�y�|�����6���9-�I������1���WD�eq.�1����&��+�NyFUU�mX����	�U�W�Ԗzlr�u��4UY�#IK�G !�e[��/q=�J�H��iW����Ąarn�D����9�e�k\���qmy��
e�ft��<�	�UQ��P�ەqL����a�sw5Q��O��t��9�}g�K�|2�e�U-�cP�'�ڐ���>����~�r�X��6��.*�zH���׮]c�����?�xr���g�m:f~vز�}�>��_㻞]��G��l�Y��|8��M�F�&�r^i����2�|F�����x|6C�kq�/��m��G/�K�.���ǰ���_��/��l����߷�gW��&T�|��mZ ��� �8�m:2�׫�E"�I#�Y�l�E�NǓI��������3@� �� G�����dv���eɤ�#�P(��W�Dmp�6�ڮ�v��8FY�p=���Z6�)C.N<v��H(�V�8�g�f�xx:*>���3������5q��?΅�G,Nϒ���	�ւ�D@�ms�VHS~�^��40(p�9PH'-JB`x��
�k�jx5�$H��[V���� �R�yӶ���E��,����R���Z�+A���y�N���� ��:2����\x��AR��3Gŕ�Y8�>�ص��ؐ�Lb^+di���<�E�*ڀ�u���H��o� �&qdox�bw���e��,%h� �2�`:��{��w�Z,�h^F����[Pȟ����1�4C�g2f	
y��EE��5��1�q�Ŷſo�n=�mY����LUcG��	��Ȭ�2��(�YQ�t�}y��r����]<	 x<ڣ�;��GRj�L Ծ����sz���3�i�p4@�i��<�/�V�%��4�s�A�ю+�=�v�����`@�S�6���	�J�SQf��|o�Z��88ne��y��Q9�:��L�%���\W�0���I$�����P�$p5�f>6~R@Vs�͜�sA�!�N�+>�������<��F�=X�^𵋋�CDQ$��cY��^|����ߴ_���4Ŕ�%߫�B�����0��Btpxx��jC^gO �V�w==�]W��͕q��_��bͿ?��Z�\ �l	�����?���+נ,�d]�AV�
����"��x� �E��4.�(���,���yT���~��O��_���ų�������a��
����g�o�r`Ea����?�r��E�N��	0_��t�B/���q��B)M&8v ����\���˅��@,�ĵX�A�n��[/���L�ݜ!M�H�H;��@�iX�d�4�D�V�A��îD��m,���)�
y�"�bqP�	
�T@PN�v����әy���f#Α���!I"��p��j��0S�w��ȗ����*S�~���r��j!2,��d�R � �(�5d�$��p��8��f�����yWG�����k�&1�<�"ڀy3�v��l�ϕk�ڲNZ#�+�.˔�A���<?v�\N&������P��ak���/�=�_@ ���NX�6rW���Vd򲜹�R����ϖ��}�X�������@� X�R��xY	f��ܸ�a�'�.�F�.��,���I�ɵ�qa�e��p�����ɼ:>>ƽ��x<�kݮ��g�/σ6.����D�9Vۍ����1ZP�<�)��9�x�<��	�JT�]��)3Y�lSD�k�0�R,����	�%V������d�ږ|�~���f��_�2+l�	.MK��򾲔E�׫�(2R���q�1 ,������-��s<$6��O{L	:�����^����:({6�9	<M_�^+��ܕ2��y�y�q؎i�+����\2�	xu`H6�c��!�`ֲM	9n%x!�T� �V��k��_jǃ�U�E��$ �}F�{��!L_#裍.//1��ٮ��m�?���	�$@��! r�ڠ���#h@���g!Nt6����O�`W̔��'�5,g��w^������k<={f�A��Yz(�qւP^����3�A����-�oϫ�|�k�"����m�>����������>����^_bpM`e���g�+l������LW.Ju��O��S?w�?���{���,�A�_���������^�dyϿ��v�	LU"��m!�@��!Ў�-1�p�����#��1�Lqv�f�{���P��rd����;@��;#�W��U�H$'��a�d"�`EE�L�D�iv�R(R�� ̬1�@�C����t+���FF��<����Kԑ��b�Qi��@�,Z� Mx���L�f�%e�8N�%�A��uK�ZY�K�lכZU�~c4�>�Q��)�m���!�����ڂ!
BG�.S/JI�FU�p�Z��p��r�{C����co[L��*�zL�k	��b���r1ATd� ن��:B����d�	<�[����a�}ҋQN4`��h�P3�ZK�h.����+L�a�s\�$�Fv��,l������N˽kY0� B�%�)\4�1E�i�߀* Ԩ�6�T�B��#ӧ��h���tL5�*%�k"�tBJO�VV���C�~'�A�����'y����d�x�5��
��]�ŋ �Iɑ-ⵔu-�5�}�^���;�IϚ�b��L0jM���@q1�H�Ѥ�k�r�q�CNv3/��Ҩ���k���ka�<�GQ�X�#t�c9^]eH���3�r��7Q��\��
��GXy^�u$��)�{�y��D"G�vz27� 	s�s'x7�n̑�q����~�l��"#�9!�cS������F�Y)��̊PF˵����E^�%�3M��\��e��+YZ	�.�6�%�U�hɨ30cl#㮐�@AQ+�),��~&�(�-a�	&h7��f�3#�`��r]�d=	$�_ׂQ:0�O�������H���E&5�2�r�n����AZ0�Q�x�L��^�&Ě5���aa3Kh��t�I0�s�R��j���(��
��lu�b����{'0�;���_�ͯb����>;��a��zӲ�	�\��NZH��q@�v�9I%�*�\ߓ&@�T���:���5�y2�2��R����r�x	
��2��V|~g�F��'�&���렴V�n��Ƈ�Ba\���W��k_��_�᜝>�>6(|��G���?������q�������9W5�Q�BU��.N��@Ϊ�tC�1�"A��E�(8���/A)���u|��XNb�]$��p��ׯ���� tQ�9q�LY�⌟�𔁴M#�Z7e3��h�����d�@��ep�pq���B���S-i*Q�%j�B�Ų0ꅜ�&�u"��f)j�_/S`��H�2��Ցѣs��^���9�	1]-���
��u�l�X���.�2��#�"#�c¬ T)��%���3$*-2��X�H�k�6k\(Nɶֆ��$�X�0��3�.�XW,�o`G�.��'Hm��hղe���B�\<�<D6
�<
{��h�5�0��lR7��q� �L�R����b$M0@[	��rу�	�:�g�EN����ўj�BG��鴷�z�V��)�AJ9�-�#��&3d�8�1tl.�P�1B?�{�Ir�L�z6��)*Kt�di�9/	Nu���}���+X,LSǶ ��`��a:-�u�����9lۅ�r��r����e�A��]�^�"NZv�e���k���L3�"���C'X�@Š�*$D��:��^_mژ��9�߶Z>ʔc��`ѱ�X�$�@ڦ&��QI��e��nd�\'@��2o�'�i-2��
U%�+UB�w��v�_-PjA�-�f��a��� (��L^;uz�܇v�q,3e���7+3��'i�8)e��\j���<c�}�a�r�R͢�g`�	S)�N(�;_��l����䒭f�2��c���d))� X$0����z�K&@L�L��c��W�-�M�4� S�E�B�f��%(�n�@�m�1�tA�#�r�N3�j6:qͼ���%���%�Z3H֙����Ȉ�r�t��G�)\̧��������~�1lc���p�z�n��81�t+s������@�;������n_��|�'�Aph	�'��3�@��B��A�h��%-�!� dR__)}L�Q�	V�_$��k�aQ�kKФ�2�#�*AR*T��qkq�ş��?���@����~�����=9�����0����я �n`�I���
��%��)NOO�aP�7_�E��.�ׁ�BD���C���O#�x��o���P�R�m��g�����cl�a0��ѳO���BD�Ո���F���B���A\�$�@K�D�lV��&#P�{�����F����d.ZM�4��-��R�]�u:K�u��[�(�(rqĵF<�)}Nt��`%oң��B���1��`��8�]mZ����}t�t��NV��m��l�eb�\
����Y��9R��&B���B2����"�뙈�O��\�qL�)��Q.�
�LW�P��Eh5�y��5%UF��$ڦIґjf�0DVLiq����LC�0�/���y���ѓ2?]�(�lE��yuu�Y"r͂GH��@���I'x2��΅����	udU	�E���GpT�2P%(�oSۦ� �1�8��b���Z��)% G�`U�X
�>l���Vt�(AY��IF�K�m�n$=<=��� �`4�qm��l����a�u2>�k�嚽� ����a�^�n#H!{K�pU,��:dd>��Q#�}l�Yi@�]��Z(�')+&S����m���J8,r��`��t�[����������#����a�*��0,Љn��uդ���kS�;Z��S�:�ت���	zd,2����Yf��$'�֒fJL)&��������b!=�!���y\W����㵋LB���%���4'�OV��`8����"O�I�S%��=_�P'��2(�`�ii�Em m
D�q*�X@IâS1A�C���Z��딌5������<�q@��y#iP��:&˨e ��9�m���	������%�p��?��bq�J��T��2�$�Fo�Ż�� �	.��7���ϙ�S�ڃ".ۃ    IDAT�%���f���^=���a�"����1y��ݢ�Q�r�H�[?�nIF&�� �	NˬКEhI�h*��;��rg�l�.��k�(��8S�A��k���e 8ؓ j�5`{/����O���^��M�=v��-�A���W�����UT{{�ṟĽW�?�+���w���>D�6�r�@Q��g)��,�Qk(�U���@��(-�'��O���1�����U\���V�y����)|��8����sKҨfͅ��d]�ئb$��	]
S(i�����ea�����T�6�i�Ӛ�8#{�^1����`�^��DR��O]K��ʱޮ����)Vf!��1�E�0�t���T!�"�6mJ�'�l��\�lRa �l)�4�*E�Q3�+ޘ�)�!2m1���f4�(p�#di-���"M���*�������),x�!,Ӈi��00�a*�1�e��i�EIpm
���A�GH�"ZR]��>Q�% �g�"�a&���Z]�,�CEGK�Ce�?:���z��
��/ﷀkC*&���0���"V���D���>������'%(�L�Jbцٮv�i�BϷ����}/D��E��Ibt!`׸�\�uz���"V�·,g,�pp��	�|���9�(�y��c8@r�EZ��V���l�$�t��b�o~�$�
��^�>�2�cTpNZ�|�Kl�W���Z�Rd��b�6�b� ��d��r�3��*	dly���eUp���%,+�r:��W�D�B7������0�,�!V[o6�m���`^��G$u�����@bq��p�q!ׅ��tE�N�i�g��n����FHMَ�v��Ұ��#el�3*�ڄH�6�tE;I�����DAf�����.p�?��`����c��9_J"<�i���8�ă����*}*�G�I3��d7ة����g�F��R�B�05�\�s\2�q��)5�e��&�[�cװ�F[��(���WLي�o2t�(aJ��6.0�-puOK.J�i�
�}�F�:`~7A<%~�A��`�-�����S� �!�Z�H��2�:�M���h�z��O�s���?��8=}�aG���n�ޑ㔟e�� ����y�B�+��h�lW�H�4�e)� IA_�k������%.�*%q!~��s)��5�Hv9��ڷ���T�������d��5aU"�X���������������F��,��Ҽ�k���N�~��xr�^{�q��O��m|��Oa2=ã'���r:��/����\\-��K�"�
��q�[N�)�l��z�������
����o��8
ct�u�ĝ��q��S�y%����� y��]�g��Z�,,@S媻�i���x�4�:�V�'O��x��[0�"K#�\xT-i&��ыD��f�c%�<6+�	R7I&��j1�4���u$���c��11��š�6#m��-�*�z�b�*�c8>\����qu9��$���^�B�w���-��R_d��J�Je�܊���\�H���^�>@7��O����!��s���ea������k��z��g�K�a&��#L.�8���5����r-��h����+����3����;�la�Ő�N[iѷ�\�𽎰8ϧu����4Y�"�qSI��Z���1iZ���TWk͢��)n�L [�h=���".N/��!g
J�С�Pg^�}&�k��A�%)��-������o�����׮�`��x�����������kCы���<q]��t�Z�(�>N���8u}����7��.*���_�7��&n���O���`�	�l�ug�)4�vQ֩z��P�*����j��J���ɦ���ͺ8��{m�0-�ԜG�����:��d���_��e�mܹ���|�U�|�4^��AR�a M;ӃM�����%�ƑariO% ��S��	��W��Rt��0��69-��t&����1[�4W�6̩�+�V��m$-J�iQ�N�p��[�S(�[o|�-|�a��>���װ7�J��r1A�C�@�1UȎG�iI�+����4�H
�.NO����3q��M�}ֹfh�;�)a�
�v�����~��Z�E�fӶ��5>x�P�	P�wt������k�A��c�����
��r���#1-��q�d���9���@����>�rv�b@O�.r��?\�����8/D�B�9Y�%������xxM�j��$}n�d��8Yc�La(]��f��~��/�~I�5��Bc�V"�f�d
Y5͂D�f),,k$i߷�x��+u�9�K��v����,+)$�H��e�HC�U!�̌@�w������{�[2�4s<v���LQ�Y;�ۏ���Lpr�ĥ��ʹ����?����_k;?�,'��o�+c8���f3w4EJ1L�=v����L�W�����Y��m�K��{��Օ���-���x��>��J�����7>���dV�-|;0F6Ĳ"p���=a�&�%���/���~��蝿��{:����w$E�們յ�N���[@�^@幤cD?&pL��j�@�P������h{��q~~&���=�o!�׌�0}ڈ�%�Im 
�d؁>.���4��3�%��kweQ�Ը$Pi��uj@T�����ũ5R�TUBٕ�'��*�lQb��J������8>�!d��k�|���uM��r���B���<�إ���{���s���l�	^y�7��`[t�6���d2��
�DH�%���!N6X�1>�]bpt��b�,�p��&�dq[tXQȖ8u�L�;�T�m	�!����4�hA��U�z��s�N��j�>�HF��y�T��iB�	�K5#���hZ���D���i�Ԃ"j�D��*s��M�c�^c���T���j�[��3\m`զ,:�mbS&x2y����Zs�ܺ>ƍ�=Q�"ƃ!�b#�:(�kBʹ`c��"Mf:�J[�R8H*��}�-a���~��7����UB~f��a!�%ZHH�O)o�^W3��fi\$�V���`1N[E����^��afa�|z�^�&}�x��S���w>�I]Ç���00p��>��B,WWXmV��'|+Р� F��X9�" ���[��]��)%"m�Y�ouZ�w�oN�$����TyS�MM˖4��S��b;]D]^�2��VZ�I�w��J���7��&αwp����g��7z6��v96H�DD��S��|h0W�-�U�����I?��`�4�p�Ɖ��ZO�VӻR@!��d�Uj慕,�]VJ��2����S^;�Ҙ
�~p ��1B��%�f�phPh
�"��LIYS-���|����Ų��b1�wOp������1Q���h��h|�A4��Y��r-�����"� r{]�:��f�S��J���b���Q�%���X�SXfWƘD�	�󙤒���=��RheZ�;؇ayR=Oˎ.[�2H5���b����`[����n"iٕ��4���Ǻ���b:���^$�3�5;;���.:�1V��T)���}6[`�C��5���[�z�~��p�c�"�4ɽ�t�˂}-�w���/=��dY��uZ#�o^]���*;��� -�A�o�_?�ײ�_̊9������g��2�7����">��/
�x��{��7	���wY
�Q)ӫK��7v@�0_<E^la�)>q���^�@����:-s5����g�x��k�{��$�p?td���)O;��"�M`D|��`��b4<Dª���]��ɻ�������X�-v��=�~Ժ�D�l�c�!.f	���1���+)&��?��(ܽu$)�*�:��z2L)��KS"qUR��@d����OgT·�����=����e��	3@�Q/�+l�@�!+!#�W���?�c�㷾�&���s?�C�U[d��y��N�8��J��E��a5|2*F�-)��z���~��}�P���[��g�� %XmZ�^�l+[uzNR�M+"��4�]��~]����1�s�V��c6�И�ײ���J�д,�6$mEs�؅i4-SӠ�܏[D󺂛?I����߄���Gjdxxy�5[l>긂U�9<�o����0Һ��b�ӧk8�5I�yv�qOaܵad9�F'�g[L�ܺ�2���t�ᐅA&��}��8�)�B9�X�L֡2���$�D��n]�Q�Y��C�@ը�<���ͦ2�����������&�R�S���������:3i����u�v�U&;�E��(�
���E?Q$��g�6�I=��\�K�&1� j?�42�`%,^J��:������	�j��5Lt�~>]�j(QM[��Z���[���4�2��|r��W-�Sa�z�!l���2�7��>�b8��{��w����>���kv9H��h@�R�z��բTF��|��7��W��5�~��_���m��w���2��r�yik#���gc.�)��J��|	(d�Xo0����
]6s6j|O
X(���5�uL���� 9����
���}�%��FX����p��H&�ea�@��aVjJA�bE�Gs�bk�pvq��Y�B�6R��?����DbQ#�l�t0��6Pǣ=	�6�����������Ʒ�A�?��x,>bGGG8;?ǝO����0�G'7ev�c������0���{�]�K��+�&�þ�7�>�0O���n�G��`V��H����0=^�z�d��XV �	D�LO�yc�!����a��[T�J����:])Y�������
G�7�8�r�,�,�bӲ����m�_w������~�?���\|lP�ۿ�o������p�����^�z��摂��p��6������0�4T	�IͰ%�U$(�-3��+\]�GQ,�����S8��YJje�\���m<zB�i�1=I�U1Y�B�/�V#"�JZ���i .�7f����WجS�F�..��Kw�m(=�P	0lP7��Z3|��-���l�nx��{�Ŧ��'3|��wE?����琥+ܾq�*[#[/��]Iu��U'�*fn�`3��I�F��9v�&��X1<��̬�`4�б��c�`�I���^^0�R`8
�ܬ�����KF�%�gKd���k}\��=��6��ɀ��ȷ1Fa״�\o`z���..�ؠ�8�����!��):�%)&���*�&dڴ�OWrG3�a�Z(l`�{�]ȟM�FpDM�fqt3q�E�ҝ��҅=R!m-4��C��(t�	�5CWr���,G[��~G{ �e�5@��Ι�ɹc�t��.�\M��.�)���m���JQ
M����J3��#��"^�����@*��nG���H��N��\ �?!����R�K7����wŹ��	R�����7O0�8O�LE*��4���Av�� ��i_"�O��=�{�qBIݱ,�|��I�0�;]�!�U�Ri� �G�:C�7df�]����������VȾ�"�`��Gm�
9o�C�m�X������X #�����`��|��mv�h�� �G�P� �#P�J��G� ̶<a�Xʱh��[��&�����2��a2K�����k���~ߗ�F���bz��a�ZgYZY���A������2��-��Ypo��ȳC���ħI,�)�p�s�����H@H!K�`�.�BRV�?$0z*��x$�/��|����8�֐�@���+�d"�!�gi������b�aO�~`#���匡r��bE�B\P�%�UjNS6u�Kt#L�[aHW�Xg�)F���}ImSs��2�l�L9����H
��5\�>Jk�۟�,>��H����H�8�X��޻A��j�D��ɹ���l��G �6��������'�*�x���1`��Y�O]�v$�̀�c�5��߂�u��Ra���F����sl�
�׹��0��C�ܸsC���>x�p|r�Œ�n7#�r��ݦzH��d��G� ,U��f��*�������=�u������W:��=~�,�A���ƿ����ί�R���p�k�OL7>��c�:����_����?�7n��;�������A׷p��>�/a�������+Eܺn�8�j�/�����m\���C<xxA'���!FG0� ��J�n�pT���
u�J��ե�n����MO2��X':�ib��ﾍ�����,/�8Bi_Ê�&�FPȦRlB�h�����6E��G�?�����ׯ�����]�,KI�Ho6v�G$���nt�,U�f��r	�`�[8<~��>�{�-l7L�g�l�3,�l�(P�ń@{:��h<���r��t'�c8:���
��J�Ơ���7P�kqt[��X��Qrg���Cy�3��t.:��b�~�'�i��J�h���`���q�n(dү�l�nʬ��D�%)?�غ(H�]�%���,�h+���>ql/�k6PWk�v�( �i���Y%�֚�fVZi@7�eڍ�����āglj�1]�A!�{���V�n���M'��7(+���b�������,��~<�`0��d�?�5T��Qm����'l�6YHa�ޒ�T^L`Y���vMGR�,6h��\�=�#�Y����믐DkiO���3��r[-����;��V��nGB������K[�VI��,2�LEg�u���x?+ �&�����LWn$���!L������H�Z�Ɉ���u��`ay3��
U����T��QJe���Y65o�'�ಧAo��J�MC`Bk�J�7�7<Gj��-�xo�o>܂�V��_g�ݝ��?��:ӄ�>��q��6�?�Go��Z���(���C�,�#Z-�w#��&�6�&E����$O��0.A�ߗ��F��^q�VU��O�~M�)�<�����iLW����� �^_X.�]��@߳q���A���l�4(`���+�Aa�l	���x{p�=���T�{A����	���]l�K�n�\S��AǗb"�R��;���&?!�ݬ1�;��z'0�]&��W����~��kb�H�}���s��~	��@�������x�|6���v��xo��cE��;�_8�ϟ>����٬��N/�y���M�_o#��}IKSF�Jmc�7D�
K��9,�#+�جe�I������ߕ���"�:NaZ�+���)J#�ɍ��ƹh�}�G���u2�gO$; ��1)(jmb�+ϳ�8	��|����r���itx�m��tO��㏽>(䞘_����_�^����׀��
�w8�w���O��� 8x�ͷ1���˟�'_���	��Λp����<��h*}������:����ʌ�7�y��c]#�kP�gJ$�wt���NW�'˨'ނM�]�شiKm=$u�[�H��Ja�w�m���1�m��|���T��Y.6��6)z�#I�� �;K�W[Fu������~���AAv��1�̢B/�LriL�[�h�T��E���"�#\;�T�����u sQO�9�,K7�e��O�����i\ �.�6�M�3�G4v���0YWa=_����Vo}vz�くQߒ6��s�&>�Z����7q�ց��KW[|�ӟA?qyz���Lc�_�pt��k��fd4c#E4M�����L�߬���-(���r�M%kP�X����<F�I�{X{6[��w���`Y�v�b�:�(r��QB*�������K/ʆ���F� q��Y����0}����g���R�|<�`�n�H�+���;>�cϦOy�DLf�F#\�ֈr������+����E����..���1��26I�%�-,�}��"fO���X�W���#\�ؘ=aKSlB�;��-\8�� ���슡ǓN��Oe��j�Xr|u� �u�+�	�����FF����'�!Sql�Q��12����D��Nz��}��\X,�s̶)����y�I10��T��l��y)c��2��
`�l)+86+<]Î��u�"ŉ܀���\��|���M)s�=�J�T1S�ܝGkb�Qv]��9�3D�Ke=	��x����y�ob�1�tp��E��ݛ7����K�T��y��ϳޒ�ѡ�p�'@X�hc�nF��H��K+u]    IDAT�VK�8с�n��ǋ�N�Ҁ0�I3����rT�؃�4-J/)��61lEP�I��fP(�d���k2Y*�hH�DM3�̶���,c��RK+�i%�*���;Q�ͦf�F��t�{�'A}9��2�У���rө����b�5{�V�wFr��iIJ�� ?�o�ǀy�ӧ[LgWx��_k�����3�ZLe-9:�@w��	����!^|�E���o�zY����)>��g�=�
>���b9�j��tvJ�	����j��{X�V��Iq|rC2�(�BA�q�\oE*@kM.�������oIP��l�]�s��ނ�0�_�۱q���?=E�닿���"Aw�����Bb�8�M�(��3�����������?��hw�OSX׵�k�������??�| ��@�a��1Y� �
����:��|z�����8���>�t{�7��F貝J$�}�%x��D�|���8<�r���>�z�<����؇o���D�M�-6i�P)���e�.W��c����[���T}�nO&�j��# &����ڸ��A F�U��e>Y�����btΦ�L����S�2�Ē����1�u	��/�[�b��#} Ya��Hq�񵻸�LQ���Y�^���h��W�i|#J��5=I,)6Nt��=�=
����-�M�8w?���9n��#��P&�⪰�x]�ݧ3YT�F����/~�S�:;�ņi�<ND�]�)�.�!���<zA �v�<�My��fאv;)$ф�H\قL3F-h��/�4�ս��~��)�v/h!�-�trp$�H4M¥���۝�ȹ(�CY.�dr���a�!j�KFپ0	f���)6�:,��}\��V9���^(�GJ��]r"�2M䆃uF�`���E������[�:�6�����To�js��iH��[���@��y� >a���hW�^h:��T3��4�&{�q{J6m�,*�.C �#v�{��s&�q%Shh� w� �h���q���D�أ4�$b�a[��='D�!h5`y"�+1|�R��P7(�~NЕ"lC��Lp>Rt'B�#�̹a�b�}4�>�w�+ZR�P�����G�6�=h/��v�q��H�Q�ur�N�K`!)���5�	��}?�$�0�/�,�-���S݃n�����D�ɸkP��(�����y����{�H`�����=�jL����Q�'`P@�B�'�f�	�	<�Z�����X9+-���J�%:�R���/�l�Gv3jA!S�tr�������e��
`I�,��k-�]�rQ�<?S��slJ�Pf�MaS�O8.�Oe;��� �[	C��{e�R9{:�-L9j��6�4��3?���"�|���o��ߐ43Awsa+�/�-�}��=aϙA����0]���}Y�x?��Y �Zx����qH=5e>�!�]�j��l���/7[�����U�W�tހ��/'�֌�C�0��y�q�
m�>}�T���/��G��E���g���k������4G�#����wt�v欥��4�r���dו��8O����������S�=�[�c2��i�گ�����PS̯.�VK�>�p�����a�5q��&ֳ����0���ŗO���~�����^�$��s���|����40_] -���	n��%zN�[�qOU7@R��M{j9r����t/�f"�� V�J�f�l)��J�E�l�a1n��m��(�-ƣ��4�~p-�s YٟV�&
8��n2`b�n"�(�,��Ə��'gg�vx$���55`K-wQ2�7ld�B�89:�|1�-�
�V���?���rA^'DZqkA2��l�FVTe2e��&Ͳ��\��|O,�9�$�)�}L'����`�WOa�d�s��q��t���"����!����m��%��>�^]
4���*jXl��-}�C,�ؚ��J;�h��@;D:c:<��&�X�p}�YjV�s��BL�����X�AdZ����.��/��g�+��V�۴/!`N�\C�+L�K9G.`��Tv�!�a��r8ؓ{Z����z���V���r��>��-i��;�_����0�p��a���!�%K�l�1�R�zG�>�ӳ��OÔF���������@���yoOZ�p<n7Ki��m��)�=���KڝL �ϝ.j�d���Җ���㖍ع@q�W�4�m��r�B�_�W�F�Xm#i��G����v��if���#�le����ݬ�ܰ��Q��Xq+�x����j���KA
�"�fcl���0f_7L_;҃��e�C�#(,�-B�F�l�3d.����M�9��;۶��YSs�'�N�3��l#Ei
q4;I���T*	����$��]I�S�n�Im'�_�e�wː�F���)�NZ2i���S��ݞG��KSqy5�I��L���OpE3I`�l���<�Ni>m�B2����H��j@�������jY,A�9�m�y7�d�zC�L�=K�-�A��#�� �I���b���y�n=t�f�U�y���n +2�_>�7�	Ls���]��;��#Xݗq��o�Ë/}Bv�a�@y�Q�˱p��]a���r7-�R�888�b������l^~��m���o��3��M*��Q���2�-i�O..EJ�����6�-r�HÐ����3��NE��B�;��� ���Q��l��� �v������ď�(����7~�\^Nq��MTu,U���T������
���$��%����[��k��?�g��1�]�ǭ>&S�w��_����_ئ��Oj�O"<�����2��~_���[7�#�^]`0`�VW��O���{��xb�Y���%����1��q<A�[�x`c�W8w-�2Ѩ�*	�Xˈ�+�VŴ[Rq�!F�L�}��
�1H�+#e�-3�a1%��w�0�&[�s�bu!N.L���];|~��	`0��T�l����D`��'��:b�<����xLI��D�����{�nG7��g��F��(�\{�����e�����]��4J�"��{���y2�@'O%:��.6�����nL���wb��!N�}��=�>z��GI�:������켮<O�K�meVey�U��h��%:P4�pFZ��5������)fbh�!�hefW��(II)z$l7���|VfVzo^f��q�ˢ8���+�nEt�Ѧ:��{�w�{��?�A��ڄ޷	ʧ\-A����Maa~�T��!1bT�ԩ�-�@��F��_G3RTS�d��G�$M��:�kt%bN>_�(���7��=g�G�}�2�7
d�|VC'e$�H�X�)0���F��,���.;�6�\ơ��6:D9�k��H��sx��$�����ۨ����+���5X�I����:�$�к5q�3˸��K��P�F��/#::����6*�J���|�6�vѠW�RF�7eV�*E)�h�a!$zJ��ٓ������Îp(&Z�j��`0$�o�����.-���BA�j+cը�#����/�+v�4�Hb���:}�2�rZ,"��Qh�l��먷������6ȑ3@�:!�������#������@�� >+�x%n���n�x~�tuZt��Y2���߃ja�V�����M"�d2�y��A��i)�Y�����C�Ȟ�l/ۖŬܷ����f ��+��.j�����Ǒ9��24X���yo���5���d�1H�`QH�h�)=|�|�Y4	���v��5�U�Ah$����L�������x�d}�-� ����p�L��"@���D���3L1�5��V:����6�/��b
3��bq|:�9�a���x2�i@0t��m�i	��[�6�S	�7�XJ��lu	r��0a+��-�s��B7��@&[��������@�j�jW:�W�^��ϐ���In�~
G�(��$�ԁ���sg1���ӽ8�g������߼�Z�8��f
�������U����߸���.Q:eA���͔ �S��Ʀ ��fx��w��%h�>�����8��Eجn�fSp��Ϭ��dEnFW5d|x��HyF0���b�`q�����?��33'+������	;����*��|W/�8�k�`{��������ǡ{���o_Gzu���2�r��_�F=�����4Ki�=Vd���+i����Ƃ�N��&�^b���0�Z�)�o���!S�k��Yp|�H �1֑�u⸬F=��{XnB�ZP7�p�y`��l��{\VK9���h��&���Tntz��x����!�����n[v_,V7��;�8��ZcZ��#�� A��<�6���6*�*��Ɣjx�5RU��6�c�?���е Reҝ����b�xbl��葓�r��0W	W�x�]�>�`c����NY6�R��hb�ӂr�6n��m������u������0����h�3G$w��"���v�-:��Ԏ��cS(j�~c	�RڽA���QB|��t�	#j����9���I���	�Mb�?��X���(1Z������Nhn\{9�AA<�v*4 ��X�5�E<�M�!��<��c�jh����1Q���Ьn�XY�f2+E9E���80?�LrEP1����U�BmU�'ăQ&���0�->�W�Aj�:�^3�}����2�y�bQ��c��OсitJy� �Pt�D}�{�RlԻ���Х��c4����v�L##n�8~���77V1;5)NN�*�2�(=x>�wt&m�x�-nv��}1�{t?��%L�lq|m1Fd,y"$Ӎ������ή�É�d
р_4�����F6�#Eߟ��z4���=#���Ց+7`���j���5$D�'9�}��)�x���Jjs�$�����{��R
z�[&�F��u��bB:�\���$φֺm�*�삣����.!��1�%�酘���1�(�0�vc�/����[�^��I�� �3�B���{�N8���\'Xp�{����{��г i�8��K�d�AJ�x��vŸf�h���9���Hw��Cy�Qp��2&#����qQ
#]k����tgF`!�U��D����n��RM��æ���`7݇�G��MC��Pi��h�1�� �?-|�d&��E\�q�3s(r��+������dDc
]�rp�i���H�8�cd�=NF������J��z��L� ࡤZ��R��{eǒׂE�t�k5�W�Vfww1?=�[7�K��]�h�]k`m��a��g#?�� ��WϡR/����/�"�ahhD�}6������J^�����$����cf�����_�)O����%���fYs������׾�/�(���)�V��t���'��;2#]���-D�.dsi1��L!����/����0�.��|N�DNE¨��4��JzC�ӣp[ ��ǉ�Z��Gd
aL�l,��I�T8&�EF�v�tJ�P�`�)�扖�Q&3h\|�ZD=�s4��f�*�1;����8B$�0��N�3�u4Ah(���A��F&W����t���h�bJ:a���iX�x�M�T����q��A�\��L�~�<���Ө�>���]���"K�L�]�6v�EU#NF�ʩ]F�*Wo.��Rn�(NH���j6��z��.��}\|����:p��!��*�5�ǂ��r9�8B}E�[�O�C!�-tM
2�22���R,�=ݬ��O�Ş>���^Q(؆W��t�zF������HC��Ml/@~�"���b�I y�\T��k�6�&��m��8�h?�ш� �.5;��MĂ^L�� �s���"w��n��=NT�5(V�������c2���W����/�p2'Fc	���>Ȣ����7atx����5��Jgq��è�k�f���D���2KǓ��#;V,�ŉ͜[��te���sl�k�{׌l�z$�����A���5���г��afz��(#1�r��m��Sg�qE�#�h�hV��Fq�ճWQ��0?��������8yl?j��,4�́>����cm��Z-vui�V���Z(!���{���nB�D�|�Bv��耒�H�H�,�6�(7;(�Z�"2z�h(��}�Q���j��
n�܄�!s�D	F2��{H��|�r]��!�}@�`Q�$������2Iכ���-�x� j�E�*�ۆ.������?�Dw5cC��BV�=b�l�.rTm�d4L'��ldF��`?�K���Q#'�f�yK���z�)�1�u��tኚá��-�_�x��];�˯�#߆b%���a��3�Ar5���<�Y��F����6:r��B�8s�M��UL�¤�Gc�rW�ҳ7�\],�W�S(�j�{�?���V����#��a���=iB<1d�6�G��;++r?�'p�(�y791'����N�������rh����P_�����^�aU�_4#��x�h�!������Y9ĩ��H��P�m,ݹ���;"��0�����k��Шe����Ꮐ���.F�G�-m�A.����H�C�	}:�=2�&h����b���w~��������?��i���w����adL��8z𵽽�t8A���(d�G�����̕���P���LsFa0�ǳL���_|��Ek6��:jXS,�Dba�ҵ�k���B��|���V����@�kw0>4�T��������G���	���ʥWQ*��pڑ�䠨�t0�lf�v�Pc�1a��ؕ�Z^ �,(#>�a��P���1��)�y�b��tB�H.T�ai,F#���A��l/Y�Hf�8���V3,�4J�ɥk�)�C%�C���r#���aVe�^&��?Dy7���x��-���w�(טb��T,:�B���+�c�χF�	�ǍF��B�1c�T���,�u4%�vG���G8�n��n�z�9�K�36���) p�Brv���j9������v�w��͠�S�E��Φѭdqb��5���r\�p؉�˄^-�!r�h$h��#���<�G�����ó�Q��12>n��k��9���8.6����h���S�^n,�j�)���{&s��tpqe��&H#��E߳��2[�&�;��f]�$������=��&a�ڍ��އ�i��ڒt=g''�Þȕ�o�Q� �czlHdS�ph:���!�ń����#�Y@|rz�%�~�YG���f����U�����r8��Z�D�#��|9W��˺��u���85 �Z6����Y��}�w�	��*�3Ǯ�Oe7����C��Ehx=��fx��5d��4Gb!KY�ѹy<~�}Q���R�j��s������b�j��WQ��qd�A���8�8�{Nd
A�G �N��Zn�MpH�]�$�_� "�Ӂ��ĂI-��~��`��Z��敢V�Q��	;�E�g�R6�@Vv��p�-r��h�ҩ�F42"Ņ��Хl��)�T�@����6�83VwV#?۸x�B�@��{�E�� .�d@�L����r�?�Ӥ3_%��|G����a�b�Hg�*��̶�p�Bb��I.;�i(�D�|��P��|O��g�#bv��aQH�
Mv�h����D��h��������I�OL7����.r��o�z)pY}���4��<�]LMfRtS��\u� ).s݈ TJ�8�VH9P�eκI��B�;��vln����#E����F*�@����#�Ńl����F����h������/1���8������4J�:&&�d���������ZXh�}ȃ[�X����$�>>�.;JE"����&M
T��`M>�1�UNӛ��y��3��Q)��j�q��B�X^�����'F�����߉t�.fg����1�����I���!��2�^�3f�Y1׸n�4f�#�J
:��m B_��\So����3��#�*�����@�]~P�ԃ~�ϗx��-��T*�r8��V�^]Y����:2>�n�x���cys3�q�ǫ��ga҇ⱡ�z�j���7�ܝ�V��t�Y?��Q������3E���u��kúގ)�C[Xx��?����~�k�s�yri�    IDAT�����*U\K�l��>y
ǎ��k)����Ϋ�7�a��*]�a1 \�v^�Yt&�������Ɔ��\�Ӧ#�!pc8B}�
=9��4KA3(<��u���șRV��
�]�h�����C㈒�n�w�.�O.[z��6'�ln7���h�L�6�=3l� Zf7r�Y��f�(NI��B��uKoCeέ�E�P������B��$Mt�v��_�R�Kp-��Z��@[3K�1��z��05p���`l�{��]A�G�Cکw�K.&yע��.C�?(�g�`�8�V��f�+T��{�8���_C�SF�b�3<�BI�p`��]�~����i��Uvo��H!���)�[���G�����Fc�����Jt�K>3��D(Er�$>��ݮ��˃�<��^��uX��ґ���ECmKaĎ�Ң��!��.�+Y��%�C>x|nD�>ɔ���>�-#�v����NZ�Df�ݏG��/�Y@�X�=�ޭ��*B����;�q��ah�.�^֗���_��Vsc��f��N�܀���܁��O��`F�ƥ��`x ������-�1	!��F%�+*f�2�L�TQ(���;؄�pGk �ª��TC�Suw���ang$�E��꓎������R*Ԟn��FO�?z��"��lǷ�n��s�\��B~�#�&&�l;aV&0u�>C��\J�L=�M����P��x���C���	��}41-���F�z��H*�@kT`�ـNzW�ڬ�^�@9���7_G������+E\��������xPn���&�ɍ���:3�ۨ�W񃗾��h��󇰰8'lԑ�I�h�v�"�����Z(n^E3wN�
��F�Q�Ο�zR���D<�����jTd�JT�89i��C�U8Z�QM�uA)l�^G�$f��р@t֏16�����Hjaڎ���.#��6�VةW�r{�0h���٥����d�)�VR� B���-�Ov�>l���}�Ͱ@fR���;q�Ӽ�n �/JWz��t�g��C��bcaH�M�Qk�6�lR�0���B�����F��B:�&�W�ɝ� 5�����A�5���a�y���
�?�����f�(&g�Qjf�ɦ��������BKu���G193�%ͥR��bՅ�M���%��w��NM����X�=�&��{9�g��G�u1L8�>5:�}d�U��E�a��w�M�S�YMnoctllP��.�//�auyE�V�o�@��B�]FGmbt8.��ba���c�;��"�I�;��k%Dvjm⴦�a��PC�#8�H#�3ԃ���_�wOOL�'���foz*��Og�[�\�������}�o~��ݺ����9��5�|�����Ld�/�L�u�ե����_.o�r�U?�n�[�����;�xi�{��M[���N��L.���Z��������YӺ�7J>?+���ڜ9~��'����R��E���K�����l��8(U��:��j�܏C�������<�d�:ڭm���Mx}�
ray��M�#��	��#������z�H��9`�ڒTB(5ݪ��pMe�+��q�7�o�H��3�f�� #��ބ�aC�d V�v�XD�f�F����-�1�B�6�i�av�a�a��}��(�a�|����s�*J�,jZ�݊vϊ���:��|НhQ�n�a��_CoeE_w��*��8�{�i[=�mf������K�4L����(��![ձ�ZD���G��:��cp<7&��`��1G-�����*2����υ;�^�х "A3f����V���>L����A���!iǖ�L���]\>�Mx�X{5x�>�k]l���\Af��v+�r�VX�
,�&�4����QX�&�d�Q�U�f���	fPł�ZKo4��[�:�6���{��@}[��ISa�e�b8j�[���uPM`�(�Dch��H7:�J70��N<�1�Z6\�pEt_�v���Q��J�`">.��#a{c;�[���hW�1����(�r����j�'�F��!K4�e��:��_��hb-����pF��V��f������W���]��f�Ba��X�E��6�WP#�	Tvn��{���p[�h��<*��u[p;�c��EC�aB�m��}3�|@����P/��ԭ��� �t��5��<\.]�n��$&��A_K���8�if���I��N'���-4�w`�Q��Fa0��b8��C�m�������v&���a�Ϋ-M����.^}���Щf`�p��@$1�t��Ʌ��"��������B^o}u�.�$׾ת��6��Ic��T�ID�`v&��{p���x7_�3���$ڇŝ�'�Z4m�`���c.��[P,ll��yK�	;z�E54x6�����]&H ������ǆ7�A$&`j���3'QvA0~y1�����۴��A�d`go�M�t���N6�NSZCf����KD�F�Bm�K���#�,B4�Y��0j$c�D��d6��.$���b���lS�0�����I:�94�#f�2J� �Z�d��Mtx=yh�h��|���{R��,ǔ���v��6Z���Ex��5�P�
N�bix��O,���.�{����Gߏ�W�q��M1Dj���&N�8�f����-N�zԻ6�x�p���&�߇no``�3�����&��?�d#1��tᡰ��;4�Y�H&7��rW����һ1�Q3ʮ��W嚬,����o��#��]�<�/�$c��ˡRHbbԎ�}�Z��2B���:��	�*elnnJ'sjjB���Ē-�ߣ��R������m��o��S#S���c)`��^�����+ك����vV~!�ٱNL����w�dk����c1��.�3i�y�J��ŷ�}�ks��W���79F.V|z���v���՝_.W
�r��:26�'�	�K�5��n+&uX׫O�Z������;����=uq�VS#-�|��o��֭Oz�C�;u�'���$G��׿~���_��?�[w?�5P���+hk�o��Z�0�8����]E*y��
�,�M.L�Qg���948,N�)vYl(���Ri`xȎ��^���*LD��V����A�-A����L�tK�����"r�<��D���E�C��j�&A�D��X *V�(R�m�Hejp'�xϣ�9zN_�+��I��)��RPNncu��j	��
��%#���9��; ��"6:���A��D~�e�]!��ك��#��ߋf�,\8w��C��Djg�fV�|���>���e#����w�ۢY!��[��n�5��H��9����D�^F,��{�O\ƩL���Q�Xp�g�0{]Ռ` ;c�ʻ\6�
8��ml��[l-_���,Q~�h�M0Y4�<�5;z���*�ӯ��Z	�3��P!��m�}TZ䀵���~�r�ؤl6��%���hݚ^_�n�J!WX���ױ�t��WaUw�~C"�X�vu3��yH�U$��þ�c��.~����C]gt<�Hb���;%�,N�s��w��'?�p؉+�_�tb�S�t�� �X0x�QD�f����-��k�Pٽ��	Lj��6�Syt���C�D������[x�o�&Oq�%��W������'�{ww޹ ����X >'��a�8�,l֒x�����PD�����*g�RD+f;8<��u�����`b�@dw6W��y�fJ�
BiB�(�cCh�*r Q57���M��*������{142�B����7P���/! z)�s���P���䱙�a3_'����g0w��5B������!\H�(�j�!���:u騥�9�;R��<#_<�"#������]�q	vk��
���� ���V*�t��v{ݾg�����"F|a������#\ukv�ٶXD�_�f�7��Q��1pW�ceg���$���=��s���6G�tu*{�0���,���kW�9�)��y�a'p`�0S�K�VS&���9�8�,�?kX
znPDj�b��Ng�g���0$��f�iz4eY$���r���G�j���V�+ w�F�����<��	���$�(��Y�b#�����=����J��ߗ�A	�����:m�4I��N��
��Y�G4�:<p�G�Sw׶Qk�Pm9����N��-���nJB��o�bn����>�lf'^{���0�v+�8o�/�*����������h���R[�.,��T*%�?M(�1�����?��R:�j�*�z��+[A�ْ���_�;����������Qk��y���[o�!X,��^��OǾ�Q�6Sh����ڭ�[�E�Z����A�.���WW��5��q7[I���J������s�������r�����>Um��C���`�U������Ϟ�L�ǳ��ǒ;[�`(r��>���;^G������bn�1��O���xS��ݩ�����I�۩�,fG��}�Y/~���g�ٝ�L���g}��߃n�w�^�f���^}:�������3;�r��8y�_|>�I�}W���T�;��O����r��q�裟$b� &��\�i�Fm]�i���t������'~�S���>w�Z�͇zˁ�7
���N�S��7#�Y��)q[:.(�ܐ��G�ݓ�Λ���F$d����̘����X���u8lnAX��A���e|��R�Fl��^:�B	�z�m�%ؼ.�*� s��p��
�2�K	�?�!�.��d�K�2�J�>�ӟ��3O`}-�����ￄ�Q�L���[@����mF�ԑ��iU0���g��B{�ŋÏ�6������翋�E���w���C�\_Z����N������Y�H<2�������"�&aemE:��hH�߉n�ך�Id��c7c|L"'<i�Ecvwc	O>v��{q��U�om�b���c��~8�~t�}�ol`jzR� Vo����ʛ������8��b��s0��E?Y�v`��(��t�"<A��]���cchT�̑�II�i��o8��SM�Y�!�#�Ja=�D�Y@����߅�P�ޡax|ðjA�&Ao��y�o~��T5/�^g�bEP1��$��mF�`��{�����_��0�f���O��#�*@m�ؾ���;+0�]t�:�g�D�M����>��;hW�:�G���]�&Ɠ）��ob2����	t�U�Y^�;2����~k7�p�ܷ�xP��q��i��~|���0�p �Oݏ��5T�x���13B#��f��{�)Mbc�6ο�m��-�st���
��]�M���(�U�����#r�����o��[_��U�8;�c��
L~bt?|�{X<4��x_��ߢ�Ѱ�L��t��?�8z�	��v�g���RH�n����)d};u�(J���$���S.d
8���x��?�@l�z���Q1�fǑaf<���JaA_[�\�u�z�^��0���'p��#0�����~/��j5�'=���0Щ#�uK�07����v��ZKCdt�ȿ�phjiw���Z��Q��\x��9�2=Ģ
&&�PzF��PBL��^4��m�����>]��6~/�((V��9��d$֔�E�p?VJ�����KQGs� ��������Kg�*j���X�ɘ�ו�PP3L@a瑰H+�6_�r��8hM}�?&Ԛ1u�R�Z<�Z���o1��(�{��]X�|Wb�7�ƗE����]��Ll�}���@��A8�R3����.c���GG>M=���Q\)�<��l��M�]X�`��n��j�v��h��E�l��>�l�z���T�Qi�c��u$�V%剅�����?Ug��Ӡ�������/,�#yOʞ/L�S�_�xݩ�%���E�X�13G�ɭm��������e�^���߷O8�N�G�-����\������XZ����4;��S�I�gr@��}3�͌b}y�L�*u�;�4f�'������|6'�&�,^9f��'���A�O?�?x��G?[*5s##'���Iv�&�tІ�6�h�m�/��7o0�Ǌ�
g�&�ib�%6,&L��\N�:T�U�M�u�I1��]k����~�^)��m�Y�����8�{M|�����js��N>�����fݞg̬bE0<�����M��V?�j���8��r)�SA�E�L~81�j�ٲ*�n�R|4���P(��9���r�������W�3�i��B�b)��r��nc���٩����j����v�,ג��z+ȃ[��@(8uy��{?���f�����f�\K$&^�c��J�K��]��*j]�Y�j�fow:&5�Yo�N���-��'.
��ޯ�Fv����iq���Qd��%����C�V��W`�Q{�`}}]�>�z���2���T-�E�t�jqZ7�����6T�Z�y`�I܊��
ҥfʢ��0R%(������_~��D�.����Ǉ^��&B���Z��`,����� N�8��֒@g������+���cj|���o���M�칷ql�0~�!�l�ᇯ��M��߇����`:č�+�<�$± 6n�k;���
�c'1|�_b��ox�۟�)Ca�<~T:�����/`ltZˉ/}��U["�{h�1NδӨ�1r��du@\He�D�m�d��4A ����x���XYZ�B����C���?`�}���+����������7�g읥	S�.l�,���zq���L��B����m�/�	G��i�S�4\&�&g1>w���"8}�1@!h���� Eo@-wD��tw�x�����ZUN�x6���I��c��-t��Xz�G��B�_��(��v�'�b�'������O z�	�ZN��58+��%�a	� ���o�������������@�^.���wR�;��m��8|�8}�i��J�y���@yq?�2u�r���ߗ�đ�A�}q��\zg�� |�i�}�fr�F�òP��m|�;�+lzsCa"V�0}�P�u��wp;K��`��~����Mn�~�V+��24�0"�g�:���ė��\����f=p� �*bc�Q^�G��^�~	ۙM�^��i,�?���O�/�����P��?ٙv8L�"Ȕ�~�P�B�BR��~�w�����
N��0������������1g'���`����˱s�lב�l#<����]<x�x���n	�?��,��~���a?B^&F�����\�CU�ń�	zh7�����C�,�z������ �CoTD�v��l�1�� 667W�ȃ'�o��i�[��f�����`*M�]4b��.X�Xᨓ��5�<t�MNy�!gD䑢 A1�c�@2�,�fD��p`7�X΀P���=��6r�M�9ǫ��Ȏ������B�QW���&�f���-9��})nh��%�b�3��|MO��6'D�*Mb4]0K��Z�S�&y�&��h`쨱dאE!;���%��@F��#�6jjGƭj�lN�z��0e�E���&AV­[����X��k�f�_l��qtDhx��	�<&\���b�!��{/��ѣ���ŷ��=�ؽs�&z�!1h������)��{�©�)�+��֤�"vs}�+K��G?�ہ�~�;X[���H��������HI$�p��A4Zm�
Eт�����='���(�=93%���_y#Qx��,槇q����q/`��X)cus���1:6�;��āς�E,6,����1%+�����<�{�����j�=�@N1��j�7n��X,]*�{��B4��l�h��3�����6[L�0i�^o��h�-ff|�L�.��}q".6���5�����^��Fs�7�l�>ͤ����n{��ʕb�Vmy�ry�ؑ�r��l��Ύ��r��n�N��O�	�0:2��U{�f�ͦ7��q]nwj��6�M��#���)�l��k���bR�ˮ#���,�/��Vu�	e�ҝ�Bv�0QpF���t�SGS�so&7��ev7��j����V�����C(<�=69����Fә�QѡPl=�o��(�c��Q��z^�^� �s]    IDAT��6�-�S��^���׾�W��v�E���|���d���Y��1=ă��pb�Z��5�Z�kK"�u:=F�}�QQN8\�:u���ȇ���A��+4�xĊ�_������񈤚��jJ����	��:����\ڂ�[��ށ����<��?�Ӏ�DOk�4_o�Ro��x$�7��Y܆�倮��&a�=��ކV+�������r$⋉���v"�M�׭���$�>�N.��b�����\N�v.�UXE!�o� &����!�f��e�ױ�����9d����z�O?��ğ����H"�bv�W���KE�.1�/�$�s���������o`'���G���iY�(.fMM,�^x�nܺ��}�8���?9��Y,��bzďD����VE���Ⱦ{q����^���2�/�B1�q��=���8��,��lN�]eaw��#��s��\�������S��.���p=�����͊���8�A�;!|��?���)4�˸��`:������0z�#� �f}��-��{��G��������u��;,Ea�k�30�d���^�/}W⥸W������d�֑�4s���N��� ���!I�N�	�����u���m�7qp!���:��8��!d�ܽ�&�6���� �0���~9�����.z�������]zI^�C���������/�9�&Ho\ı�!,N�XV�83k(Z��el��8z���֭����36�V������`d8�+�/`qߌt2�Ӡ"��D��A���ÃG����g���)������&�;T����d=�H܏��^G6�,N�p��y�ø��;x���x��idRi�3[���i�PD6IP��Wn|K�^�$>���!����[taߜ��(�v����wQc�d�	�ߎ�k�ju:|���/ �ZG��W���X	�`��c���7,h���A-�5�V�.prS��4z=t���+0/�O=��>��=A!���S��r�Ǯ�
�.#����z��ד���/�.ԙ�g�"�ߓ1��FB���@�4��×�f���&t1�r�s�&]ȳh9"&*I�n��(8v��
�ŧLg&�}�f�6Zm��	N]�Ux=d�6��-O~��yC�)�F)
�d&:p���{"/�S�Q�PP�4���.�D�و bڍǋt�R���3Y��$Oq�ki-�­�
M'w����i4z^��E�Tˈq�oi2B�A������h�'f���3bw�捱�Q��qܹsw�Rh1��f� fX���;x��9������}rX^�-�/>�5���2)2TY��-�?��,ӣ�py=����ZS�@\��6"�����p���ܯ�LQ�ż�����L�M�T.
�cm����#̝ם,������ē�a߾}l0�=O_�)�~�=Y�˼w=l�q��%N�=�����Mf�Y�X���A�<���n�k���b�����b��O��r�Qcʮ)�U��I�"�g(�M��k��za5� Ԁ��G,���i>��l�nO���$�k@��Y�٤b|b�R�)$R���Y�SH�o >����5��?/񙚙|a�rz$�Z)�U+��w�ݩ�u��p��2����/���8�m��N^2b=p9�Q���Kj����`���!KR�Ĭ:��/yV{t�;���U8��0�>�p��Ha������گY�-IUh�8]	X�S�z�Q*�p��A�rY�,^ԪM����(����׶ӛ�9v��i�
TLO��ܪ��R:��bf4�~��v��x�J��b�'$7��E�f�f��w7e��Pzvb�y�}�5̰9��������א�lahr�p��(�fa��8rxmS�}��3%�-k��\���W_$$N@�'��B����$����޼������w�����'�*���;/cr!�bہ��Q��pw3�ˍKo�������@��+@�z�Ch�������rZ��ۈ��C�^����x���N�6X$Jr�  �"�+y�]�����0��Ի��[oIw�ڍ���D�396���Z}�<�$���/ �م]����E�����a��Y��N���G�������a��x�h�^�V��i�p�ZE�8>�Rs�ν�^ӎ3����\�s������8��]x��KX�\�M0�H7����"zJ�c#(��c(4���N@3հu�5�zy�,�uaV�p����7��j����w��x��w��׿��7�����>�Tp���9����p��e�����Ԥ���v���iT�ot=���B�ْ�S_����X�H�44sKp�k��ܶ����_������Ep쐘���î��p����,����mc{�M\{��1q�'19�jׄ�/����K�hUXz5��� ���3�����>t�Q�{�2~��/|�w7��b4>'r���&��|�$ng�Ѹ/��e�*[p��� �/܃��u8��cc(����j�$��3�I*X_��͕s�'��;�я��n��՗~�'9�~��,<(�K��\������[�q�Mds���[�b��=�;��|�,..bq� �F�P+��8��iU%O���Z���+�ˬ��s[�����Z�V��f�*�=vI��[ĭ�$*-��b�*d��ۻ�S��1K��Io����'�R]�v*+�����D�'�9b�Ȇ��l�s�wQN�c��M�� �4b�=~�q��CM��׏b�-��l� v�&ǉQ��V%C�lC]��n�8���>f�s�L7 �5�U�>[�8E�R,���c���h���l�M��y�H���"�#�[�9�YŤa(P��¿G� &Q�<H0E�C	H1���������LI���Ōn���n��jߘ�(fjk�R�����Pn��*����!G�n���g1:{o^�
W��}g�L�`zb�7��{=��ܾ�h{}�?���.Ȃ��u<���R4����8{�,ff��|��e)�X �9s��ξ����	���nh�P�U�2�����te�C1�Tk5�|L^�K��ݵLLO`��2��~�ss�0�
���ۛIY������t���S'y�B^�����3;��񸝨�*x�]�c$1$FO��̳��>���3���3q2ş��{�F�l_>kI�;~���K�����d�&?Fgr�$Q�f�����D�jVP.�`�͂�r; ф!�0��R���m0���N.��f�Z���d�v@�ÖZG8@%W@$�A��E0�)h����*��*¾��C��w;uhz�K��&:m�"��N�v��"�ӏZ�g���;W�Y���E$<$zfr.;=�1��u�<�h�]�|�|�m������o�L?�8�'.
?�����h��V[C��.W.w�Ɏh�ga��r�Ш��wŐ�U���c|<���i1c���Nn�N$br�"�+�:��E`�`�5�Z17����f MV����`�������*����}�q���H�&�PlA8�$�z7o�¡7ű<����K��(沸q�58�m8=G��|��"v+l����o�艣T��O�/�^��F��ۊ��x��1������.F�a�V�8��{��^Fr�:J�u�{Nd���&đ�����˗e�M�
�9�G��ċ���1���<���05;��;KRl�N�8ܼ�x��i:q;d��뷰�z�<�8>��p��ul�l������9Q����S�z�i?r�4��n��{�����P��J>���i���y���LO��o~SNd�������7�8GdȄt�2V��¤�15q|�gp��e����"�qܾ�"9��f�B������*N�?�!���:��Qd�)��]tZY�~����}�зy�R�`���>��}�e���eL�p�p���(w9jT0��?��x��`rj�ZC�	�x[[�F=����C³l6[��'>�P���Y�}��6��Ȯ�!\���a��*&ٲW.���?�K(u��pAo4���h�3XYYEph��[�U�mexkw���6�0�����ᥗ��k�_�V��h:�>/�.��C��f�2U��Bl�I�x�4���_�5�� �=�#���Qd�2�1��X�y��tNw�ɫ(V@����$���~�u<�سx��B�P�����̼Z"�r�67Wq����m�J���3��_�ܗaS�8~�������rI�nF��)�а���������m?x�)ܾ����~�~���(���Qo'N
��P��/╗���/��鷱u�2�w�	���Z��<���u�p8=(ժ�{���������@����P�����a'S���0ឣ��-��L��@���@�ϫȢ��E!�{�4|�U�c������Y�L����v��*	!����U!����O~��L:2�1A�0��B��|��J�!n���i�G�����ad��0f��(��u~wc�Md��F��=�[�6Ьs4mC�U�ѣ�p��fl��g~� 7������|�{�p:���k�L�������l�<�k��qq�7[-轖��� gxBCk��T��fp���Xݬ�̣?��� ֒;p�H�(W�8��.�u	�V��.���tj��rh4�X\�'E��ր}�Uw�nI��I��|�,o�;��>��DG���߃]��W����=�$I�����Ҕ�����x?�~����#aC�)�J�I����E�r<�D�I�'$Ḱ\`=�~w̎i��{���Uu��C�_�vb0;]�U�_~��>�c����ڵkb"��uckG��l�
y�q�B"w�W_/�X���x��'�Fp��q���^�ԣ�tF ��W/#�N"_,��~@�6��H�Va���1�f(H�{}Ǐ-B;8���}���	Y�I��a��X�9��B�8���-z�0Y��'Ґ6jDŝf���g�����R "��|Ν^S�i��D���B�A���#���\n�X�F�n��׃Z��\f�rQ�.\a����a8	2�����ixl�-q��X���_�J��
r�F�)�m�������������XVW,�rSi�uhj
n% �� 9�f����E"���R*�A&����5%*O�zg��;���_�F�y�h��.
��՟�m���� e��*`��2|(WP��-�'��Y�ꊋ��T��CvjF��LNT�$��~vĖ��^]_A
K�~/<܀�=�a,/N��n�&�p8��U���b�v͡!��rn�P�vk�����cw�����w:��C�օa(�J&��q�� ��0��H�?��K����u����h���o������̱���9l����7Qغ�q������P�������+4��2&��g��o×Z�q3I�Xߐ�.�ɢ{�����7����Ϣi��w���m���Y>����uYX?!h;)2��,9�}�(-k �=F5��l4�k��;j_�p��%��x����˯]b�92$�"`:Ck���ںx�;M�ㅗn@�&��q��9�b�J�*�2��bb~]o�"�bu�M�J%�>� ��|7W+�*��c��4�}1����Ѳ�Ėx�����>���[��%�lkЁ��`sw^�B:�Fܫ 4���Q�+Al;�V�b��c���O����B�`_x����	(�8�L�zq���x��g�'1Q�y��ۤy�)|����i����+h��P�1��V`5�������]������=�Í���df��Ц��_�o2��/='d�z��cg�����A�(�[��S����ڭbn�$6��P���^~�A�z�˅Tr�H�2���7��w}���gp�U������#x�=����MY���h� ڍ2�Y<�����߅�Ct�._�����Z	�~����O���3!�D�hɚ�)���)��z������9��&�*�|�}�_<��|�i�R�8u��R�cI"Q4�u�0r�T��=�
%t�[��^A�����<>����GϽ���=��o�"�8z�1����qH��Y�Ԫu�zU�Z�?�7h�6p祻��_��z����}x]&z�&lz�)�g�h�-����t��O���)��4U�&nn4gd�X���<7���(�A�L&Xd��gB�mO�;��C1��5�{���w8F��m�L��q����0(J(��9��0a�Uʰ���[N������|��a�@�`>yZ�/B5Np"����ٴ�1�R�e���:E�c�M4���"�c�
���n���A���:7G*ũP&C��6IQ�tZR�v1�3��E�ę�0���!�z"����\�=����2�s����w�VeX����{����)��ƹ�74�ӄX/������Yᕊ�x����N��/�%F�Mf��G�����bAH.!#A���X���,b�>�NT*�p��)1�稙E�T6+����Z�	�SռBˠ�i��@
K����8s�Μ;�g��jO��)�RY�c~<x�t�%��M'�����lN��j�*��<�ȱ=��8y��&Ǽf���F���o�}@��5�uL�N���CĔ�$�q~�ۍ#�x�n��"�:��j��it��i�O��i�h�Nt��T�x4��KΘ�<B^����o`h�c�f��A��t*�hxV
�rm�I.��^[��\�n��S!�+{�9��۷M���]*\�!Z���	�,c�X������,���DᐲΩ5:��4G贐�J�.�W�lLO���~�N��0��R��D�i/� �׈�6�K�,����-�7̢�1={�O��ٯ����.
��_�WF�ƿV�* *��':����PUS��Vf�A��y�,�W�/� �GE�1�V��PA �VC��^�T0H<�a*G$�Mń���୕-��a��%�����fL`�ZpOT���R����E��F*�,<:��探ӛ�6�}a	7^�k��o���}�c�رQ�������*��`HP!xT��G6���.�[+"���;x�Ca�|6��,-�C3_��˯"���SWP��pe� -5����8���^T���h���AY<�� |�ڭBZ僒�R���ǎ��t�00��V����(=��:����aAɁnãQ�� �HaafYogϟ���.���b�{jy�(��J0���p�}�bs��+׷�ȣ���	Q�;��8|�&���.J�+h�v��v�W���&��}x��_��ɷ����O}�c0�C}^���l��Ƥ�-V��e��&�
��;�a6��3k�3��ޙV���x �a!��(k렍���/�KDsw��g^�������.����0���!n޺�>�,ܪ.n���lCD8���,���u[�F�����tH����=��&��F�m��c,����>�X�0���pPl 6{	�6�yJ�^+���֨b�P���E,���e`�����T]E21�t�8V��U��p5�����&>I	���|�݂C�������c��}�޿���Ng����ă�B�tD2mu-,Ea,C�`?��� (a<n!N���-�
=���c������5����S��ohdL��̊�qo?z�	ă:�*�S����>�W_����������Qi4pP*�}���9N����������;D�oⳟ�U���ҋo��?��Ȥs�U��mTJ�C��[�$��������kh���{�_�T֯`��_#�5���a�@*�D�TDP�A�w2��kЕhA�=B�ߕj��a4�n�u�k�JQht�������,&��Ӱ�j����ÒE�s��Ս�XGA�=L�D����C%�tvVx_�;�b<|���]"[Exiz��a%�	K,c$�LT��2)���DQ�E���,�_��u�mx�)��ѠЄ��z�iL�pxp,�-���YE�?���������:x�����I�&�����\�*_Ma�)`��b��r��J�A�s1<���U�Pu7�h    IDATm0�0�:3�]
t��^��D$�no K�a�(���p�+��9�g��
�&h\�]��1�}8y�$2�(.^:#i[v�k�賾�&���+W�Hq������g�yF
Sr�X,
��e�Ĝ�y�JI
���������<|>]���{�>X�%��MI�
�����`/����µ���԰��7�(6q�t~�D�'�M8Fs� ^~�A����Ɖ@s�Mt�?�g�c�cj|���07��ٳ� 6���x����A{�����������l���^xu��o�����L����M׎K��ɡ"����z��Ao,|�N��N�&��,�A[��l�#��c�������\N�8�t�1U�)v[���y�:����{��z�@҈ؤ��=���*��bQ�{�d@��
oR�(p$�˫D*��^�R\C��-DCs��LQ�G��L�Z�Hx�"�"�۶�&��M,��pin�1ƞ \J�����Ŏ�m|���'~�_���kI
���a���1cD
�S�/�9P0��N2�T�K��8���@̬�K�M�E����"��5!mP�s
�y<�!��\�G�X�܅5֡��b,J�۱�3i�� ��tz#�!(�F�4��T�h�?�1+h���5̧u�<E�\�KT��]H/�O,�o>�-ح
���,�=/�{vD$-�;h���L�(쾂wޗ�ґi�=����a��>�������΅���Q�وp���2��;*�U�{���΢A���ح��1�Q��������TMs�� Iq��ڐ{Е�_=�D\���z�����t\8{�h �j^8Y�=`TX4�CS'�@^\��Cx����W�č�m|�3��h
�ۇ��@@���4_H���
��������$��u��c|�S��o}�5̟<�dvZ�Z�v33i����ҙ��x������b��Ń��D�u�I�w{Hd����D����t��)*�jg�zkEO�#��"Z���~M�����V7p����ħ��������_����F'���F:�.��%ܸvG���\����g�g���0q����`�k���aw���:�I�O�B&1{�p+q��䷱���`�8�:�Xʵn�[�HF"P�9A�U�#�2�Ž菘@0�X�4������ڍ��6V�%TF=��25��A�w�|�A�̧͒�?���_(�p$)M`$�k�C˅f��hЏ���l��T�1Ώ�<�+��ݯC��wޅJ�-��a&5���}A�책j� kk�!�3a�L����x���7��=\�|�G������Όo�X��z[+נjM��]d�g�ɟ�ylm����>#YɅbM:sll�dj5�s@~C
�NJ(�70�x�<~�CE������]1�D�赚�Y�1r��Т�(�+�9�pRh����c쉠ڠ%7r�׮��b�V�a�ȣ���S2�����c�(t�BrT�8�A�((���i� ���`<�_��?;h��4{�F��ظP�+E&fE�1x�Z ��>�����0��AG�Q��ƒ�@�'�Bͫ����V�`�|N�8Q>�T�.�*8z�4�'�Yr��!/�V[r�ÊK�z�mT�%��p0�n��iA�X0I�qix��u*��K��� �L���DY��ժ�{mj���,EƠ�G�+�a"��}��~,�}KE���~:;��_{��gΜÑ�yY�[7��p��6J������kX���H�Nt�j^"mlƋłܟ�奿��ln�����ƪDE..͋Wn.7�T*#�3w�u�P�X\��d�x��w�z����_�zU�x<&t�+o^Q����H%��@�"5�I9V>^��	ϐ�/:}69���8�����[[���墐��O��cH���Rԅ#	G=N#��8FRī�P,C��m��Y�D�˿sJ��my�3w(�ԀF?2�R�t���E+Arټ�5�E�[u�HҔ	��0tw�h��>ʵ�C>B~���b	vo�d"���m�@G�9��/L˳6��a{�j�ݦ��Ŋ�	�@P�q*w�[�~G^���/�C���$��� ÃN��>���^5�|�!�8���� �w��i�#����g��n ?�� �))&��\>���~ᓮ�R�mԄo?���o�򿴺+���gC�;��)$چ� ���>hJ��X�n� �����,Nԉ"���T͏��:��ҾI f�5M[��8R�������M�胛R:±\qMǸ�G��X�	����Z#�l�ȞDb��,*��H6���x��o���w!@�hzx	���n���V�e�0ҧ�ҸP)��H���(�S+�Z=�S'Ә�S�\A�����k#<��H.���6�<�r3����ȸ���"����#��`��Q�0RB�Aম{���n��(�az�b)�h7��\�J��0��6����zpwv�wB>����'���t�^	��iX&��+HO'������~�7p��ø��x������� �{T�,s���F�����6���[�N�"�����Kw��}i�@V�xzy����1�������r�9�(��1�1;���m��s0{e��kP�j���\��M�]?�)����1}����+�q��g
�Pra~�,�,�}��$�x⛸r�&<�_|�@K��X$ے��]$�q!�����S�e=��TK���JHGU�?9�fw��>���T���s���	ϰk����S,��&���!�1I���sQ�:v�������S)c8Y��1��qmgk�m��Z���� zܘILϞ@�6��v^oS�c�n'.�D��\�ܐ��XXG��:F�}�_�L.,M��9t�6v�n"�� !��E�� ?Fė��Wz��~%_����5���Hd�Ocw��^�B2��LnQ,3Xly�
���k{=�{�hն��<�ba~#[��+�8z�|�8��[݇f��G�ըcH��F~R�Һ�Ǐ�O㑻�ۨA1��4e{ԇ��O�d�.�{�#M�G��6E�^�-��)4�� �e8D�x �:��m��Y�����|�ל���c'���8��Š��Xb^������bh�m�L[����������S1t�L�9qu��H�%,`C�
gl��$�n�Q,D�8�^߀����̆���4��A�ʾ����&ǎ�PПPѼ����-?�8�A�����Sl�/�"w�g��
�����5m@�0Q��vk�f'N���ڦL;�/�BWm�
K��Yt�dg�,w�fH�jJ^g�v���$�yЁ�g�H-"��B�F[��Dڑ��h�Z��o�<�,��pJ
o�cV�\Y�3��jӔ���E!����9�(�[�����2�S�Z��h3�H>v�|��ZYFԤ3P@��*
@x�2�U���8y4�w>|7&�_��Wp��I��E��!��6�g��^m6���mn�M���F�R�yn*���kx�c� ���B��f�s�O�>��Lg'���)9QQ60��ޟ�吉4�#h�!��	��n2�t�~���w����.�LL�k����F�ۖg��N�P�XRƵ��Z�6�[��
w�KE�Q�����=��Y��xl��H�R�}��\A�ӐB8�Hbg�$���sg��u�{��u\@zr��.���Ea[C�Qڶ�ru��G�����b��f�B��p��DIG�X�NrGiN��tJ�1�����.K(lۍn_]����H<~�[��E�SO��������^)BS#�J�:7�~��(
{��#a�c�Fұ4e���CU7��
;�UI��ἃ�(	d'�a�)|X��:��n�>2e؇k�G���9rcՇ�7����F��8����~����h܇7^~�_�/<pG� �p��<� �l������CFR"���O�qk�
6�W��{&�b�6��� ����f��i�GU)�SG%=��/��ڊK�S�)��t���0���25&ɒe'/�В�4Ȧ�*7=+�Nv�<d�Uk5�h8�ѽ.)Z;�D��{~�-��'��Op��Y��_�,�gBhR��k����X۸�o�H< V?}S�#}gO?���}���kx��O���l�<|F����P��c�tv��wN!�C��q����\�h!��ȤxÐ�d^'r��ڝ
�PϿ��0�sD0���Hd�_YA��G@�c}��vv0per�|$|q<��� ���������~�������Q��#���y�嗿�ko�3�`(.�Y�Zt�| ����%�������>���++7P��)l5v���Ih8sb�2�[�����q��hW��Sȣ�gť�jZ�����3�0��X��sG2H��(�K@|ss��.b�����]CbZC�]��Բ��o?�h<=����[8r�*�>Zm��M���>��8{��}x�a�$Dn]6@���/����ia~6��}�Z$��ؘ�dp��9���.�$p�:(Qy^E�pa�����[0u�L�ΡP�J����sX�;��~�h��I,�.�|����k�V��D��V��wG8�A���t��:Ś�#��4\$�[�t���<����m̤B���Q�6�U�]�u7h�Ʉ7{�D��.�96b��t���3G��D�	Ǫ.����N�>�`�� �_X�1��J���u�mif�p��u}�#ccF~��T��`���gk�/ݼL,��PO�L�r��e$��ca)h����J%��K0�I(#[���E�B�b�^��]�7�`f�)���H"Q�`��i�@��	��(�,f�ră�Š�r�;Gú(�m9G��8�r�V)qw&<�0���խ=TMdsӈ����Ph.ߧ�!s}�7�F�g�����ꫯ S�Zks���[Mt5i@U5�fko �xj
�d�����+�����H�S��D�g��x�Q)�B�6�K�_�o����ޅ��c34y~q���9V��Л���D!_x�y)�h2��w��[r}U�!�t��<)SD�|:�\K(l��{>m��/�B�(���l�vG�]6>-�cmm�p�t�f]�m�;24T?vt�^���	��^)�� W��3JdԙNQ�2v=E���$6U�*����Q�S��k��#���%�y>r-�{ff���Z���eb�p�^�]�VezZ�_쁦RK8w�������:��3R`ѣ�k�[k�7���$�T[��Kf���{�2��\�!(#�E���Z=�=w�4
��I�}�}��P�֝"v4�u�+�P"�>y�C���4���,J�bɄL�A'�ѫ�%��[B"���L��Ng #x�ٹ�vP�zæ5�8{�}�����m%ϼ��������_�]Em�*�M	�G��hl���ۓ]n���ҎD�6��I��`4qƚ\�BT>��y��9sѿ�_$�rSB*mt*�Tx����0�	��b�Zv���<�7._jt�6�6z�,��K�� ���Gl��՛/������8�LT �G00��.���=�S��=⨋��a5��xse�԰���r�]9�+bn;�C��@d&�B��a�{��1k8F�!�|�"#�V���.^@����~C�� N`l���O�x<*\
�� v�3�P�x�����uy�*�<���M,g�F28r���S�-�SO����[,�2� v3�]50��x",���s�b:w�R�V������&0�FhT�b{@Qh�ä|`��g���� ��1�g�f���
l�1�����\m�����]t
x�G_Ǒ� �y�))�N��ΝZ�Ȁ�e`k�xaZ�J*�X"�4#�.�J�"��K�������/ j��3���(�A?z����Z�S\�G�v��H����<w��%V<��3v	'�x4�0?-9�����{���k/~;��S3"�Ԯ9Df~����}!�&����y4Y�54{#�N���N{o���h����#1vrc�hx�����x��ҙ,\�k�\(�Fx�_�G>�k�k�Ǜ�+(3n2C�]�gl`�+�K���Y߂��G��0KE$G�n��ɳƣRX(�11ě��U�&u���J�=t;U��Jԕ���1,�ށPp���1	�"G/��T*;h4�(�7�PISk��=����J�G%UA����Ă��24m�Vc��*4��ٔ��Z��rR(�`"Q ����o^c]�0�x�1�({T������>űH`̠�7e�	�=8�����Aɟ��o?)o#(���r2>B�T9p��2q����=����ǈ�n�iq�	)��8�.R��~��49����$ۚ�olDY�8�Sđ�f_��ӄ����sw�FD���Bc܋��k��p �猲Ue"�^,*�U���V���ߏ\&-<�S{�BoȞoF��T����]�!��ۨ�:Z����~���v�������=�����W�. _�$L`�R���s��Ɖ�9l28�ty��5�Ba߲@#��ȝx���4�"Q�C�8�#B~n��wQl�H1�ރ4���ٔ5�=�Q�˞MRR쇶D��סM�h�z[�N�Hci>������������(f�X��Vz�z}���	"�B�OӉ����d���b�����V0v�Z��i6,��~��!�/��?I;�m���d�E�
EmA�5U��\C��w��XX�d��p��i�4+bW���ws2c��`��K�L�Χ�:��8�,ŏx��[[&{V�B���Ws���XoK�i ��83���!G�%b!N�،)zX�����G���B�t������9FX6�|�]�"�']�7O�4{Gu�fNl��"�LI�4̑p���i�&=��pR10��c���.��3��������/�����z�uZ�\	G�=�b<vb�f^e���|h�b`-�;h2����K�9�bU�`��@�*I��!Cs�9�"Yմ�P1��.�� �Nc1��בˆ��"U�vɃ@Q#h�^�r������4ߎ#�X����ކ�iö���������q<p�G�~k���ҩ�2�1�y;��4CU��M��c+�-�z��Ш̶D��t%�ib��t��V	��<�cX[��g�Sb��7_��O"�����4�����6�n@���~9���Jަ��Z��f_�%�����a�DLzu}E^�{�[$�m���*hQħ���]�!��F�����K��j嵻���t#u J��4�J~�����(�'h�g��jD�F3���8�C�����W0q������u�e�u5�{^��(�� �=z�{0���xd���C� ����G���ri��A"
�&�fg$5H��V�g��:�}��i$�1��~LO�G��cؾy���Ьo��7����v��u��~;^H�z�62��$��$ӷ�>&`;�p� 7��S	��q�7�u|���;?�A���YF�sI|h7k�˫���R���թ���©9�4��~,^�"�y���s����������aLF�Y-�Ef4��Q�0���p"����ć������	��%ٯ������S��+7_�_���^YE25�O�$��*�Q.< �h?M�m~U�w�A�(2��]\߾���F���6���R�,��)F��_�6Dx8� �}�������m^��*#�D�4��p� ��]s��9lu%�h(� Oa�ʥ�P�2�t<t�F���ٽ�K��U����IvϠ�7a��=p��R���b,��Cܒ���j���L\v���^��o�9��� ���
M�8<l�o�����@Qr�)d�a����l���:]�x��{6T�32f��O����#��DBx�EN>+����Z'^4�`L{��3=J���:{�NO�A��.�X� �� ����/,@i��5ԡ��L�$U���Xi��G8�6;m�Gf�S#NR��L 9���-�gQtjux=\3:��:\���jՆM!�����1��c��=E�    IDAT�jß=��7��vy�g%]b<��l�?��'�U��,
����씌��Q��<�Y`s�~��iY�k[�=DUo����S�z��R�q��~'Qd{k2e����ŦiH�BD�ga�t ���� }��*�G�O�X��8:�����!T+|�Ͽ�P$���K�`wOF�,wv7�F���G8{�X���V�����{q��������T��X�p�*ED�]2���K̦;My�|�L�%s|��΂���2V'2��"�����u�������A(,�T���^�$-�H^�S[���XC�܀��o���tJ�n����
R�*�"|�Z-�"1�3Rd�p����s���5r!����h8(�q����� /�7c�Ǐ���"�h�W�c{g�*�s*u���	*�Ƀ��aG�_U������7H3H-n\�����{���u�������?��ϻ\�����6R���~���o���)��!+s6�cA#:ק�2u��a��|b2�H�==���p{|�u���.[�ݒ9LSJ���p�&�"�}���>�m�(�
N�f�v��^�l"���&|Ѱ��
yy` �a8�a�J�����֎����[�Lb��iاZ ��~���I/>��O��3�[_�^|��y����g�6��\�G�N^(�W?|���&���������Źsǐ	F��157��2p�#�x�(�U�x���zC�����
J��F�o��O����N�yPx�LOD����7!�ք���87+r]*�H�l���3^���^l ZG�=���ag�2��>|C�:��3hY�{-���X�Z��O�?���"��2r����F��=B�e�PE�������B"�²ţ2�L�N`0I���M|���_�4~*�z"�+lb�X�ϯ«��UT5	z���n��ud�I��(�r�iɟ5�=\��8\�`ku�+O!���׮��<�j���ܮ!"C�04��0e�I��ݚz�� f!��)7p���#�J�x�\�yt�>���V/�o�!�\yg�.cv:�v����};}QlZ�*Z�<�IJ�c���H4�c�?	w(���U�x�[���ܼW#���
6����k���?�odJ�N�j�͗�{�U�8q���rS��0���G*����5<�����؀�6`���(@����wÂ��dM�ⱍ0c�4R��r�حn��,��,�8W�8���2�B)��^D���ʄc���bQC�Q�p�����u����ފ��Oc�x��Ex�%�^g/"''U����q1�-��a&��qg�u y,�|x��	j�<���Zu��Y���eQ���
����{}���xU��h��#�Ns�c8�0,�i_◱dr6�S�0���Ðq��a���(�7�!��.�]d�σ��%G�B����(<%��B
�h��o&R%�m�h��1=�hW�"��0-J��k��F���.��C1ZOg�q����L&!���}M�7��
y~}h74�BLNԮ.}csI�q"G�+'c�p�H����dzr��=zPC����@֧����T"&��J����Bςpw�����Cv6�dz���v���h�i��3�?�o�_����(;f­N�)B"	�q�=�drBg�Q""|��p�w;ߘ�+�N㥗_�E���`�YD��_��4�l�y/�_��H!F �\�>�)�������ގ1Lv�z�:�&�	�,���h761���=V��3?F����;Q�����[�G�p��:T�N�#��G�l��{����NL��v`��_F����*@��Z����wǻ�׋�0~�L���w��'�~S�/]��s���ES����$���4���Y��E�=�>�g��snw�V��P��d"��1�tk�*0�x,� ��V^�N'h�帘��Z��clٷ1b^i)�6�.�0LD�LW�F!_D��� ���dCV�TDA��}X�XA2�$Q������6��4C�*�2O��l;�nG���x��v������ɞy����\�x��U������U ^|�֪^�/��B�ۄ?����ob�CA�00ىj�&�#��C<u7^1|��0}�r\�����c<tAS4`�w���͝�F�@�E٪#�1b)��T[uc�z$
���"�m(خk���'�:��ÿ�c���ҝ��&�4�Zv��{/Έ���xםR��ٟ��;Wpra3�e�-7�1��p����]TAm�#���¥��Uv�ѱ�P�|�c<i�q��}�� ����a}{�.^B<A�`[#�4W���).ر�Y�h��@�w���U(ȃG?4�����b��bz�k�c�p�
�UB<��D|Z�0�A��)4	�eX�%�����*n��#�n��|EK��Ex���.�P���gv��Q_�/>�m�v.�F&�P�R��'����N��(�tK^���Ht�0tk7d�
xT$�a����e������|7�O���GPlmKa�G�G�${�,o"���J����"*�
|A��^�/B�z�r`����!��n>s���[}��1I�a�нBW�0"�4HTK����CB69��HĿ������p����w����������c�)�����7��16'8u���� ��z��H�j��QP\ց�=�ހ���.^�rK
�l�M7jm>�������� 9�Jf�{ 6�r�*���6�z�"�v���"a�V*���p��=�x���@����Y��ܽY�@o�@�[A�S����n��Lf����jQ�g�~B:1�X��c�a���!��+yA0� �ZB6w	��,ڕ���}a&�.�)�p����tʇfg���Ҽ�����p�Z�j*t7lcx��yt��9�C���i%a|̢�-�	��L&�L0�{���ʾ`)p�x�QILsg*eɍV�����[�s�x�qDH`�&_љ Kn�{�@B�}���j@�
E�i�i�c@��@L�}Zq)y�г���3��aFt�k�
P���
��)���B�l*�!��7� �����Ex�c�DCwP(��4��z�P�c��%��ŭU�y������!mp�``;����D� 6us��@�a�� ���Dg����(�� F���e�V�F�g"�F�U�r@�Ir�q�:���p�;߅�'���5�u���2B�3�s�����X4����r�%Rq9�X�E#I,9�v�t��=����,t��Y�����3fhSɯ�ȓ�xI�F]x�<�|^M�'��D�
bob��3���e�H�_�Dv-4$�@��\G<���an.�V}�k��7��7�Pl��a�P�.��Iy�V�e,--��Z��5���r�:r�b�l�	��,�W���X���=�l�sq
��2�i6�±�k����;q��C�L��Z���$G��26&xѥ�ť��Y�8;Z������W�Ӹ�������<굊˅$
{�Mҫ0���\��A�Y\�����&�� �`��l 6A4�B4�1֓�}
�8u��r����9'�w��I�,P,���^F�g݈�/����G�x|��ץ��tZUuT�>0Abj�ܼ���;�(�^�t�А�E*���~�z�`���	<nū�'��xR���:z���܇��#{���m#�/<���I����+ZG\�}�8�	��!�7�O�hk ��0�A�#,�H���� z}�
��&\	���"�d�&��ғ�\��ɦ�(fs�0��A��>��>���u�>���Q��x��K;��}�9����	t�����Tx�.�;7����Oc����τ��o�>�u|��G0��׃�Z�x��ʂ�z�"����
�**Ɠ>�"@*�B�N`��Hs|7bSs�r��K��3�N����Ə^~	_��Ęk��e�����y�����=-�z�Z��H����jc�G+��dav�,�͊ׄ�,C��Ƀ��a��\ƃH��j���HH�P���G07�ę#K'Q��Jy����xl��X��el%d󘟝B�:D"v>]�+����c������]���bc06��ib����07�O<�z�,)z5r�g\nML%��ٻ���6�1?���6�����r��kװ�K!� ��0;�F��#��=��?�����n{��hT;b���:�I�n��<N-���lk��J'��x0�FRpdb�C����@4�E��G,B"��l�Fo�h:�z.W��0�\88X����n����i<���t���٬ �ȢبI�U�����\��O�)��2��o`y�(�vW��
b�ܮ&ܬ�h�����7��Xj#��Cs`���^�Kb쎡�U��,�����D�|s�@r�n>����_��0:��(}DBz�T��%����{Qm�2~�hF��=*,"M�̑�׮��֠�Re�K��Q��1�8}�"ҳGe��B��n����AoC��^��v�bn&ŶDiب�0�p��� Vo�1���H9�� ��7�ZD�jhvWpP�.��l:�;�N#��fa�^yQ�n7z+{y�C��,��b��EX���53z�5�{��`g�LdlȈ��!�o1����.i�݊؃� D�c(ND�U=��D��_G����cn)�h�?�۫H1���[�ښ�E�?�9"��cD�:�U�=d�LԐ�FK�����Z������IK&���ƅ�1w駀�Y���m�����a����
_����aj=l�_��.!�S��hZMb<��t�c9ۃj-��;�ࣟ�$0����o�	-ga.�t6o4.��t*���U�^�Tc�d(�3l�G.4�	��H!��A���&Vn������-�kz�ɂ�	6Pt*�vA��|F�D�x�2	X���9���G�R[�+�.6��w�|R��iX�RUs�Q��]��7�f��5��ea�)�O��f3Ϣ�h8��d:-띜���6f�q\8{B�ൕ[����	&0���jqM���,�z�yLBA��KX�;*EVj*)�FP	!	� ��壋��o�g���b{m����<r/f����'��	�Ht4���o��JG�nң�@�NCo�K��V��/�P;|[��Y ���`-��u�9#��C���=���;�|�8��;ⷨyuL\��N���w���]LFM�*��=8�����=x�1���G���ʵk��f����ZY��(� �m:�İ�U�TlF��N'��m�ձĢ�#qll����nbi��)�eo�����tn��K��(Ea:3�41�tib"�N��aj�(��ֱz�GHģ�B,1#N���=FF���3�* �����ݱ�bjP�!ͬ����},>{������?���l����#�DX��D%cYm�(88��s����-�/�8}�	�<���YgF&g!��E�Ʊ��!�M��r$�t�'w̃�׍�d�T
�b��V���2�cm������~�w�K]����?œ��>�O�n� �i!e�Ŵ�υ��gq�w����~�/���X�$prꘈf��<����	�ͫ+��w�W:@�k"7�ð]�k�E �!u!�.g��sP�`������0��G�_}�;'�/٭7Q�ۆ���̧?���~��_�$K㟙II�^sB��AW�Q	v��BQ���w>\4^�d�����M�{�&f	'�gQ����1vp��K��&���xB`�`H�9苧�+om!=����E�
{���%a��������r�gƢ�#Xr/��*�;���,y�$�)���c��a���OA�P�QK>��Ș�����[��2��n�Bq�����D.���Ǒ���F�5l��Dl!�P,	�Ff�N$��i�][��檠zŃ����"hH$�Z��\zYx�4�epP-:�:s$�֞i��y�:rd���hL^�Gqc���n'o�̙w!;wF�g��M<��?���K<C�J����>���S�\��͛7����@,D�`O|����_���������%t6�������KF�"ZFz�c�����I�n��R������W`)qT��������<�4��s��s����H�IJ�h*X��a�Scϸfƻ;밳.���+{ʲdeɒ(�"�,� A �����9}r�i�y��co�O�F8����y�羯�?�{�����`�Y��*c4��Χ_d�\��wo>C.�B<���aUq�Xg4����:3�P?�RQE���X6��L%�f2BM[%��#��R,1��B�ڥ/4N��~ꍮ2����D:��i�3Z���l�b1V�\���������~�Ç�ࠔ*3��O���ڨ��T��_t>�<�;o�����28��Ox�9	I,���5v��6�z�\S8�.Z�*CvCcȆ/p��f����:5���|֢�l�Y+�}A�4T�\:tb�w[�;&��2tն�:�?#�|!q+N��a�O���u���IS+zK����nK\2����� �h�!�$bC)Hu:���x�`ԇ .zh���΍8�t�4��S����f�;�y��ټ��4�ʙj�J�D�Z-��&m��B1i�b�+b�8)�[$�yn,���i1X�X�v��[�������V�8����Ѩf8|xF4��al/��vn=C!��p����.:15��B����Ti�j}�"�V3��H=�tNiG�V#R-�B�=�S�NYO��'���2	H��\��:>Z��`�����բ�E�Ӆ�ޓq����D2��a�]���*ܹj���/,�5K��8�e�"��b�����Ã��n�ܼ��ԥ/�dl(��i)h�n?Ŗ��� �fV���������Na��#�Ci��r��0+9���V�l*��=��j�GO}�?�A�_J�۽�5B2ʗɔբ�v��&��O��mq�w[�C-k�,p"_��e+E��~^*����Ó�5�������DA�I��m��9p`��λm�6��������l�q��EF�dhP��Hd��Oh�a�n�I%���X:zt�*��C�?���!tV?O��y��=��a4���Fg,����dpx���v�79{�>���{��CޞC}}��Ϩ��b�H�?@9�Q�C��Lh0���<���:W~�C�a��:�@�j�J%2rX/Wp��j�酸�� ) �N�e����Sg~����?��/�^~�w~?�x��Ͷ��<9��dC���61E ۤ����V�ǚ=���ELfek�I�AW��,�I��
*�9�J�>����ץ.�NSK�V�=&-��R���Ћ���s�26c���ĪN>����R+�3/��W��u�A�ZF���?�J��C�|i�>�(>��./�/�ȕW���a]}�kt����4*FO��+�s�,������S����$����'�sK��� ���Z'�'x?����D���]N���l*������̓O>���7��w��#Z��ˋ�]tGr�T�%2j��IuddL��- �O�2
�Y.JG��"�t�$���Y��]�e�;ɨ���D=)ƇB��e���md�{��%�=��:"Hw�m�FWiw��'����Pϭڬ���aq�S�F�����vj9{��V��S�����ehX��˺U�+��kU���uH�P��筛�0�T�kA���&.���P����6��=u�ȴ2X\��>����?���q��V���c'����y�B0Hl���4-��C#���l�q���S.C������Mv�~�� ѭ��!j��v�l9I&W��>�g���Vd����o��w/231�v$���!4Z�:�(f��!�^2J.E�+cw���g�����.]�#EʥU���z/�Ƥ3R�}ר�2��t[$�u.��F$o�_�?88�({�2e��U�ԛ&�~�_7h6"���w�K,��%��ޅ�vM��~��Q&&�D��5�H1�S��xW8����ZEt�$��R�EG��3B���ș�R��ɬ@��f�=��Ԑ.��T2��1
�=
%����Hp䐒/�n%����Ԛb�1���nG�dt'[R���D>�Ι��̏�Q˦�����܈�bt���r�i��\    IDAT�K����	�Rj���� �|K �Vdv�ֵ��l
���;2� ��u�+�������ץ�+�胅�*�	����b9qJ�������I:vc�r�DCLg&��|wke�F�ҕ����J���G���K�
@���Q�FS�''n�t��+�v�7��h��v�K(����y\G?I9���ו0��L��c�����l$7X�u	M-Nة�R��5W�VYK���Shz���%1}��C
3�7[���cd�9�}�e�_��Y���|��*#�G�ߠ���Г.�1����N�"]��N��݊Jj�F���:2Uf{P�Rt���#�@�ܤ�#�:1E�A�?܇��V�q��RG��"N�3Y<^�B��&5:���*%D�$���a�Z"�h��4�;�4;u���� �����GL�*}ƨefF�	L�.&���6e�KH6nWO��>*];�@�j~���~����ZBt&f�����=���k��^/�O�����;���2o\~�_��'9x��dV��E�U�*����{,�?A��jU��S��w�� ��Pu;]�켧w�E�-&uP�J3��c�tj�,?'�8�E�#�\_ �Q���"�x���㊃���/2$��p�|&�8�rm�'�)ҖH��z��>��%�Кt�9p�,FG?_��Wi	5b(����&����-�n]x?{�M^z�iΜ8����j���C�VS������4o�~�T,�Ph�j�D:���� n�S#LM�#�������!����!�1�ڔ�J&��FCEkTڗNu��)��D&���d���>b�~�U���������L��K�^ItjL�i#�=U���RI�^�V:!ѕ�hI>L��l��طo�v�L4r�F��b���Uu�d<��C��M&�V��P��f��S�#d����sӘ�U�ro5T����Z�s�����ם��#��nJ�7��S�vH��[�G�1�h�]d4�Wϥ�m��g~���c��_��w^灓�X�،�ŒB<�K"��*C�P�ao]�x)ǃ>����z�-rh�O.��&��q{�J�lcp�(���\�����EU{\��{��[��U4&��+w����J�,�TYx�{15.��V4"��J �r�Il���SۣU���?��f����aem������X��&*�����Q@�J(�%����`����n�HW_cs#K�5A($]�V�z���b#{�h�jYX��ͭUY�����if�*�-ŖAud� 9�r��]*C�j5�]'4 ߢ��C�.���TFg��Ǚc��&vpK,� p�ױ���e/��>�c�,K�I��w_�l407w ���Vt�W/��Ç1:8���I^��3ln�V�VA��`�Ѫ�t�d��'YY�14��3L��W���p�uܻw�����8�>�O>�F/�Ϩ��k���H4�S7|�^��tb5Xiu�$�{8��.`���'�#��j���V.b�ܡ^[��Pi�Tף]o�1j4�5��|��`+Seu��,.��v������v�������~�o}��0�*ahss�ё ;[�;Ή��o�����G��j�Hx��,�Z7Wn����ŕ����ٌ�4���:E��Dou+6�tܑEZ֌b���	��o����;��f�z�J�����"�i@Y�8lv!��B(Ul:�ɴp���;�uZ����ٱ�t��<�����T��Zɔ�tjz�Oc�X��&[Wia{n�.z)�:��跁�DxIwO�R����m��5{�l��S���
�uBch�CqtPZ�ZӻC�$�&�y������)�@q���ت����"�D��x�
���*>��Z�>X�B��t����^b"�e��S��B��A���jq�,���X�2������۷�����v�{zH��J1�F��d7n�go����;y�M#�����o��@�[�������<r�j���'�_u��{�\z�i2�e����x�|����6:}���ޫ'�O�iu�h]%oS���V�d�|�����l���:��h/JC6��1	m�2NHq"��x<M�&Q�v���u?�?��3Y��&1���pk:5����<yj���J�O�q��1izf�F���T��Oom�)��h�e�/.[�\�+���5���8<�{��` d48�7��]�Ã���Z�Q�_�}�U�纼~�-��i��ڊ� X�V!�uR��9~�(�N�����P�F���%F�*�j��cI�U�,�rI#���]>O�a��*�a&�U��*�G�%�Ϩ�[�2�V��N/����:i8I�費�'���N:��T�j�B84���bq�4�:c}�q��Pcts��cJ�����U�N�;D:����8����:n�f� ��y�h�Z���TϹ���;�do�z�w���`�E(l�,zkM�dNmN�����kW.Y�09xP���f���Ӵ:M�%��RÕw.�v������v��<�2y
��V]MUe$���3�z�B�B�@����������_�(|�����l����i�(a���$$m�L��"��?�dwiw�����^���3�n%�ge�:��=:�8t�ʌ�tz؉D��{b޲Xm��1+��ePz�vC2�k���m�E!��)}���[m.�+�"��O?J�i����'�}���h.�>}��ڽ7y�G_�`(3�o�FKˉ����I��hWK��go7�xG�p�rj�-_.b�YC.�F:�M$������C��Q�f�r�9�Sj4X���U�r��N`����d}���Ť�7=�3���/���029CGkDk0����2�/�M~쉈qD�b�Yo)�� i��(��Lk��0�0�246N�X�ș�(=֝��&�\�n0����,��m�zզ5ZU�� =E/V������]��&��|yG-*���l$cI�&y��+�y	9�T�y�-�ta|���S(]�n��^�,�
�j��@���6ÃnbW��يmq�3#���x�b&A�Tb|j�����x҂�>�?�K\�r����m��"��cؼn߽�;o�̓��25��S���K��B�������y���\��������l����:v?�s��8\�7����V�����wjm3�����3���������E8�O�6��S�v֕�iuQ=��E�� �����𞳟���i��_�.>�6^{�Ze�˪��--wt��n0tU����6�.��6}̞����RJ� #xq���9աVJ���6����d�K�U�i:UD�Csg\��DuJ��i7Yh�0-�k#�`y�.?y��<|�!b�5ں&V��jZ����x�>xB���@���kP���ʱx�5|"��ث%�����g�ń=8N�TV�T&CW\\�KUQ0c2��ܸ�ä��iP�T�w����9�?��]�G]�.����6�Z�UG���PU�#X	��;-���]e(,�|�#��[S��z�m#:Akk*=E��T�D��Tm��ִ%<��_�=�D��PwW�W���FmS�f����kur�
z��P��\6��uu��*׫N*˶��卯�T*�Έ&�Z��Iu}�~r�&��C=F�b��~��~�3���kJ6�REAM7Gj�*�o�H�"�:���ٳ V����UR�/����o���fv��o��h��t4m�,\�[��Kl:ɯN��>����Sb[K�,:�:u}�Z����D��^��B��=�^�����)�C����duwz�"�I%�Hj�}�F�* F�7養�r/..�*h�	H��&q�:�XV����KgQ��r�B�Zc����SIZ�
��������[+�h��jv��\(*��Er����uE���*.E�dM�Z4�a�O�e��ۄ\n,��v����D���x�N��aq��S/�V�8Y[K��RO��Ѓ�q��q^x�T��O�f'��~J����z�R�����K��DJ�X��F]��?�!���{,z@a,�5/-),��6�Uu��! )=r�y<n�u�Ɩ�W�������b{e�R!KS��E5�q8�px�DR����n����vv�h�z��S�+���B�>πB卍���'.�_}c��x���%�!���&j�?@����U�_��z�i�nv�d1U�D�����W)8F��[�^`�������l#������R)���1�Td{�
.a$vZ��<>��ɮK��W���@o�hB�Q��eA
�\�P����7|��Պ·^����N��S����. [�Xu�*i��uc���w���@���P��e!K3�4�p��]_����r��҉-�#C!������9T��BShu�*�.;���1:�^$�S�͞�7�J�r�������6񺖾��,,o1��>Ξ���O��jYE��w�������*���g��x�d"�����Y����������=�OO�&iU�����$[BS��K>��:�z[�ݛU��i�zs��X�љ��:z�#s^.�������Ḿ���de5�V$�78F2SA���r���TѤ��rb��8�����(9��~C��K��+x�NM���K�����)&���x&�?�;��Et-�b�09�*l�i���:p��
3)�щ�&K��s�c2���]��D[��\I)ǣ��v#ۼ}�2�������8� �J_p��L6?�XFm�~�[���cS:�z-�v�7o��Bc-�J�ѩQ���]���ɦvi����0:���R%��9�q�>�+\|�.�^y�S�N1>��ѩi�n�P.�����䬺2_���r�(�3h�y����Gz������*G�߃�5���3�����5t��w	�[�m��/��2<<����(ڏ��7D�V�7uH������WW�bwXU����+����u����'���}�P����o��<�'�43�xm�35�dIH�{�@�*�0�B���HB��܇�<�z"C`�_q�]d��q��U���So>�љ�N��}ܾ���3@�`�h���>�g|�k��>�!��bgg���b7z�n;��X`h���ꢐk���Co����e�b4aw;���Em�2�]�s�K�E�z����ԑͻ��N����#�3w�4�dA-�b��'D�Tgka�Tl�Vu��D����<�;�-�CF��4C� G��QN��0��;\d�	4�V�QIۡ"�����(�Z�f��t8�ΆQ���Jg�ёΥ�ZS�PVb��[8-�k�3;�T֚h��%E�H6�۸+�+qbKRk��\�m֫80)��������N�`�W=�)d��]T�F
�v������0!md1v�8S��&�۪�F����L��/4Mpl�d����6���G�p�PN�r�&2�h94�w�|[
'�=Gh���v�9\|�9v�����'~�ɭ���e,oh�-n�W�O.������!|N7�?���8��V��R#�2��w%�D0i�^�L��SFm�&�j\��٬^Օ����úH'k/�P2%Պ��E����j�F����W�"��IŬ�QR���(c�D��Ba5�N�`J���կ�V#kɡn���-�Λ���H��b�]F��g$ɫ:hҁ��)ʲq���G��f	���|�݂�^�$��v)f�����d�	�mKFJ�5RTJ�Vg���fPX����iks��=��O�G"]!�������d#�)���#�w5T+�:CoT�n6��V)�D�$�vqu�P�>�(��^Eډ�^�"(�f]�G"gP�Ma�œiW\�[�vZ�jy����KLM�S�T��#x\z��<�"��0s��`��ڳ�T:ʹ�SJ586EGd�
F�M����-2��{�44ܺ�¡��~�Rja�9�Q��~��� n���T���C���j�E��~�������"U�1=3�(b*m�j�Z[x��>/]��Z]��଺�v7;�@Ĩ�O�E�R�z/fP9�F���f�o��C_�W+
_{���(�����ZZ��j[�C5�=t�.*U��j\�0�`��0�U*�*���_~��#�)�c�U�pHZ�96V���0��t���{wA�x�V�f1����<ֶ71���Z%�Wq8�oJ�f�����6����o�qOq��lEj��k�I<�o������+�y;��*�}�|���[*y�G'8r�.��K�d�%Z����'1K����_�����\����@����S,�B޷��d�%�-�CQ�5�U�P�ɧ�x�!�%a�y��9�\�����xG�UzY��*�5�;���F�����Dg&����ܸ��6�|d��H�d�ms�O(!���՟�ld������rwa��#uzr�-�n?t|D�X\��s��C�q,�>4�F���U���T����x�]*�a�C9/o�L��<��3�
`�Ł�.��:ݎ������ec#��Nj	���.��SG8xl��ś���N��k;m�-՘�gc,�$�����|��_�������������p{������W�����6I��C (̻~�?�I�g����}��C�c���s��Cg��n��N�R.��k�o����`~��_��1F/^J��FǄ�&��M�uꪐsY�������ҕɥv	�����l��~�b�<>�\��Z*�FL	#ѓ�R��e�N,Wót[�ވ��12s��ƀ��P�Gy�Ur�4V��[W^`o�u�C:N�"i�0Ś�����O�Ѹi���i&����h���*�Bl��<�e��w8>�"ൡ�����R ]���/�.�r�_�w�I�.ڒ�Q��?���kN�`�H���gD����}�
��V�9��i�s_F��RM�vv�ދ��K���|^�#G������}��A�Z����y���x���!��
�|�P��$bIH��J4iZAqU��Pg�驤Ӫd�����:��R�t����!����)Ӝ �e���Z�T�J����K�i��fG+E��Nפ�lYKw0�-Tkb{9,���b9A��czb�R6O���phuR�I^���J�'�G
E�S��%ZZm��@*]$����8|�,��{�9����<J��F�����Qi>[;kJ�c���ʛyR�;u�O}��a���O�X��x�w.���޸đ��s��O���$���U�U-K�eq�2��o]���^������
Qd�6�7�8]fje9LȨ]�WN:bvg����Bi��b�Z��d4��#��Q�4��l�P�����~;�n�|������0O�ա�@EP�Z%8'�A�Q6�����p2��Dg�b��]e�������	�K�N�X�2}�A���(�=%Wk4��c�����CC<^$_7�:���a4�f��T$Υ˯�������웞�w��02�Odg�R����f``��LSSa'����$����ݠ/�ӿ�F�g��ǈ�%	�Chuz�����h\q��;�)~.Rg�j����V�g@1�i����*�=9��iB��u*�X�nw[U4z1`�vI�H�,+ٴ�Q�P-l����Ѕb;���~� �D#��t�x}�au��xMɮ�!
�:���@��`�064JY6�~���hmT�-�2�К�[\ ��������}���l����0�|�����^es�evvĐ�At;2bPa��r��}4JQo�����0�b�ѧKN_��!=X5)����@�F��o�v�^�i��b��F�l��������?땕�]k�R*f��Lo�n�d^L%.��c�ZE��0�MP)Z��o��S��yur���Wʼ��L��	���n����N�/.ǎ���m���P>}N+���з�$%Ж�Z�΍Z�?�T�F����V�~��#ln퐌up0<8O`h���]����u����0hs$N��'ϼ���@,�Ũwa�;X�����5}��޺H�o���A
�$�7�`7h��qfV��;D��߯��<��O،���E�QK������//�2:<���b/�'�S��#��"�M<�V#a)��#p\9��\0-��q��t6�ſ�&�ڣ�,�5�x���­�uF�a|���쵷�d�з��L:�<��j��a� �V�ǒ4(�c"����!~�w�z� ���,�`�N�]���c�l    IDAT�no����P-�avҋI�Ak�Q�:���2:u��o���A��%!�%j9T�^����OK�&�ic�'y��Y2Ֆ2��L�/�`vj\	ȷ���.�l���*Q#�{?���i���g)�K��o�������Jn��j�~��7��Y���m��$9r�g�=���i޾|��ϱ�t�9���5e�1�-hE\%*`��b:���-�_�!�f��a�ԧ�I��)�e�pK�W��OFmOT���FK�Y��՟�������S���CF���Sߦ�������S�dЇY/ё5>�Z%��A�ef`�~�Cǩ�����)�L�O��wiQ��&&&Tg�֭�dgj���n��mrd�N!���c���b���
����$ˢ6R�e���J���W �V��+�|�|�&G�T*9Bc������z�L����>����j�*#�h���7�����v�j~�l��yT�H���� �.�gO���ݥ;dDW&F4W�r����c0d#��:����O)G���\n���%���b|�������4KW/G���uЩK޸��B2���d���%b�D[�T�:) $�I��@�P�iH�lDKdk]թ�Ua( f]��K��䔹K����fI��ФEG/���L�;ME!��Q�<r��%;\��B[c��0??���C�-��N6p�[$.e�YT�F�O���Dw�z]
�m�٩7ᅗn��h��~{���£l���|���Wn��Id�6��B%G1�b4�[�dnL�C����'X�V�S�#�u�nݾ˃�~���ҕbWۄVEd/��2�m��.��o��&<�>�O�}��yS>B��:f/��*MG�a�,���*N�<N2Ʉ�����$��ҢV�����0��2~u�����ݛ4�bvJQ��p�]X,Vlv�:h;ݞ���(@�*G�#�ٍq��)��I1%#j�׏Ug���jd)����mU���%/=�F�Z����Ũ�B����R]�J�H$\�x�ÁSTMIA�������I���'������?��q���J�1���UQ��֚�*��n���+���wx�'9r��A���RL�4T��=0���K��	�ל�JgP4�F�:d�_��&��8%JQ:���(��EL��˵.�����Ozœ�]����d��S�<�:�zM;µkٿ�V������&^�n�|�m�4�3�n����w,#�Z+�Q/.�&N�8�z�l����Q�A;�JI���"�PM��
^F0; �=3��@l�S+�5��ww$P�!�&�RȋMx�r��$ck��E�2���@�RIi��%x-�\3r��Ja(��ށ�ݒ�`��Zժ�Z�?����V^|�W��ZZ�C�����=���x�d��nBt.n�'c�XT�[��V��V��j&�q��a�W�z}��XY��nN�n��`��Y����揝"��c/c`ď�]���$��]��PH�'Ze��4Q��O��L��������
־A�ƦI$�,��%`?��;�t6�>?C��>�}���;Y&��MF���'�b��ݻ�,�]ejl���n'ဆ����VL���6���rcT3�;PF�L��{}�յ-^x����]���j[�m6��Mv�6��T���Ơ7+¿�(�0����KU��V6�]m"w��U��C�)M�ܐr��yQ(���{�&�j�Hd�������X�F����#�ts������Kb�h��c=����R���fnfDGΝ�0����O~�����?����m�"��uZ�ވ��XX�E!�č׿�}�*j���?��O��_�1��~�鉃J�-Y��i�S+d0�m�V�y��oQ�-�Ȭq���|[h����Ko�[Q
�f����P�C���es��G	���?x||��Ǚ?v��XN��<>7���V"ģ��6��,e��k�<��Os��c�3n_~����c���az�2K���Q/�Ԩ��K/���*��rr�2y����!7��cg/��U!$���b�ۨ)�H�Y�lf��{o���9�z���GO���?������b��sc�1����e,6���T����9ɭ�(o�}�B����W2�T2�������!#Oϯ,^�c�0�0�,����;��z���	WpWx��FR[��KY5�+d��䰶���*�a��Q�?z�z���+�8�C�C��&r��a<A/�\SÂ��$[g{�2��*s�^��&���'Z�$cS'��3�č��)-�t�\v�F��n�v-I��İ��������O|�ŝr�;ܼ���&#�~:�&��'���Ӵto�oh����˰��KWS�R�樐P���4�qC���t�F��$Q����ص%4�:M�g���Oc�^�(lF�":��Y/S�`�;���j��^F+NIJ�x��:�GN�1Z�z�M�o���H����b��(J��z�t�M_à����-���+7�t&�ؼru�-������2�;��9½���a�l���V�Dd�ѡ�BeE��\8w�6À7E���<���>�
Z���s�,߽%�k�O���duu�[7.�����`?w���hQ�F�v�'8p��ӳ��G�"�ߦ�)Ѭe�V�L˻gA`�F�rj{�Vj�8V��s���Bz��6&�g9s�9��Qy��[Be�0;�_�F<^+7o�I(�gltR���!104����͋��{���#�M����*s��՞��s��ϳ��Űd17��2Yl���ʈ_�$�R����.s��;X,�V�)�q���a��0�i��J�'�=:'V���,��HjrX4J��h���ok3Y���aqY�b�4�YV��t.��:�Ւjmrl��~��<�����r����;6L� ��q=���Q\��}�f�%hIQ'-)��]�'���ʙMbR�H���;h���P�Ѻ2�H��r�kT��<ڝ�:pIG]iz�hm���q�g��;��;F�R�+V��n}�Z��2^L�t�=��R��[�c�"��$�|��0ݪ�5�1څ�i!�/ Q{��&]E%�HPmjо+尛{�IK�è�V:����\�v��.�{�$��:�b��N:���k�Ŋ$����A�Y��38j�,:����A̤���J�fK�n�R������F����_�)|�'���Z��2s�J���v�i�U~m��PY�!�WEޕ��������Э�� �#�a��4f�Me1
�g��/�����Z偐����Z���A2;1�F)5B\7���\oR�*�dQqHk�1�i,7X�cx&YZ�(H��#��&��'�����]lv=�B�S���V?��|�}s�h6uܺq���6T؍V�}��`v�qㆊ���%��6�n$84�biu��c����?��W�z�%Zո�l��:Z�� f���nZ��5�2��ѯF��{+��^�5ٍƕnH�F�!��,Pr#	!_F 2�,:����*
s��28h�5U�0aԕ�Xz��B�ŉ0�����GO+8�3 Q[UV�x�[w/�L�>�)y�#�}���[fp`LE�u�V�_4�D'�Id7�E�1�
�^�F�:���I��;�r����1�^��j��ʋ5;-$3{D6V�u�%t�M���]��\x�\,Bd�2�R�P�C�X���.�B��B�֡k��>M����_�.^���=��5��r���=����ki��k5g�k2����q���9r�d�1�|�kܻ}���?�Y.��l�nr����'��jL�k蔖8>&���m�.V�nV�����lV�]q>V؋�R�`:,F޺v�;��pXj�y��=��0���]A���/�mn�2�#،m�aF}�I+�W0嶹��<��!�c����x�[�o080���%7�l���y}s���I��h��4��d1Ra{��j�g4�XN24R��R�Z��r��Q\�43��ڜ'����^��v�����(]��ǎPL�X��Ma�N<�E1��G�bj�N l�x��U#��쪱��h�,:*�0�P�������YMQH�á3��&��a=��X�w�������YcmC�g�X$JJ����t��F����n�$��NWi��e�U�)BAD���,�[C6O:��1ar`/ӡ&��K;O-��Y+I]����P��u�TwO�\eT)�M��Ӯ��h�۩*�f"�������z;�s���51ҏ��n�����n�Hu$%Hl�3�*�*�[�%���H�؍֨5�j� �t$S-��YV�;,lW�vsQqHG���"]W���F����T�06�i��>�e&+�ggY�}�Օ��g0�ܼ~�.����������/�{�c<$�*;N�ܾ~~�Rk�T�e��m������(� ��:�ؠQϣ���y�I䍤2���ԩ3�*���.�hL]7U�q��-�'3���*)�ɸ��� /����U5U�B�C����^�:�SF�F�����p�,�z�� ��:�D�������Μ!��^�o���[85VnwJ*����
�E�E� �W�q��J���ŗ~F`d��H�X�����9{��D�bN���9s�)�bk|�_ef�>LzaO@I����=p��)������(��Lt:=ݷ���d��B����FU5.����KdHydO�����m��#�����{�$���H,�c���*�0�2��Ƌ�������mICk��W7�z�R1\��ȗ����l��@�mZ�Z��J @�j���:�V����:�	�^��V'�	��$6�䎛ɗE/?F�\�a먤*M��R�R�7$!�tD_���}ӌ�-��U�N=�JSeo��b��h�=�S�k���}�i��	 �F[	X�4�2)�*a���-�	�6����:l�/�3��ބ��~�����?iU���&��͹��m��0�\�h#�.������Xk�����U���_1rD�9��{��+m��a#]�1{`N�M��W9>��a,�.IK�E�����[jr�Q-�	_4`R5��e�Rl�Y\ߢXi�nh0�CԌ�󾏣�yy���YY�C1�����5���V���J{ �����C�1��~�z��rz�����S�ZM�h���^"��fTh�-�ʸ}.��v���S!VV7�w�}������~�e��:V����2?�$��ϫybG4�6�N�KKln�)��ͻ��)(�
Q�<�Y��X:�
�P�+a�,j�t[�XW�D$�Ct:�q��,3����M�s��oar�9z�Q���g����Y"]����@WUa�5
����<F��驃���v��F���(Xr1�P�l8�D�RO%�I���߻�����* ����l4ݬ�aht^�ؽn;z�*�<4�ҩQ�䩖�
A_}c9���~<.?���+�\d�g�#��;�,��q��6��d+%:+�B����:x��������<D:!�V'Kk���;��������H'W��������9p�aB��؍n���c�:s?ӳg��)����_�Q�(Y��e`d�L�+�_�N_���ӿLb��KO_edh�Q��7.�����5�"��Id��=6#���`���դ�n��G?�'�K_�KZ��
]�nK�j�<p�a�N�9|+����C�D����n�W.�����Ņ۬�m�-�+��W�K��Xq;hYB�ϏQ)�0��IU��^̐o��L�N$�zq�A��Z�E�&�.+�^M��!ٗ��o��_�N�b���V��j�FKp#�+�~�N�x��an]�i�թ!ܿ��|����J���Mv�J�ӿ��dc��;4e��(G�]�t؜��WIŷ�y�kL�ˆ^���ߠap��L�z���~�]t�i���VT��P-�:vv7͆d�K��u��`T�8��9���w��{�Y��M��B%��Ǣ���#_H*xp�YSzD��L���e1��P)cr8�����.�	^��q{���OQ�I�j��Q<n��K��������W���&�ȸ,j�}��_�Z[}�S�2I�n�:�J����qC~PA[�]��m��quM]�v���Q��,vC��N�c�O�@�D���?�8ξ��\��r�ewg�{w�)���j�ՅU2��^���S�qo�G�<\8?ŀ��[\�C���m<���Y߼�7`'SH+�g.���T��MaD�@W��,ӭI!5�F���?�$gϞ�d���[�����X����	� �BO�V�l\�UK)��N�T@���$�Q����! �^l�	�诳�����l0�)�qz=�i�6���Q/��jy�>���N��HWE�Uq�L��_F�V����	�F�)�Jf4<q�o�`p�����(C�A޹~��^��!�+�2 �[e5�^����������8}�ׯ\�����yjt݌p�����O|Fu�l��ۡ)+�V� �l��Th�ҷ4j5���JT��|&����Z�Y����^��N�#��;
@]�����`,2 �+㊰��k�h����$Y\|�`ȇ���@O�(��u�`_F��]��dP�+1u5�Z%wA_��^�h(b?Bݏ�5�pz�v[�V��nm�R~�r5�b�;���p�P/�R#��tҔ�)�&1{Z�хF���*6��b&�E_������A���yߧs�yr��ٜno��^ �@ $@�<���,�&]�h����Tٔ,�%ʊE$A�$��p��y�6��0y�g��s�ݮ���t��j/��L������y>O�*^���A�t76s�N���؋��7yQ�&Z�i:�Y�B��J�.�!��m��)�+���|�omRx�_�_:��`�*�C�x�\8�"W���?��/v�$��M���byi���Y9��{W���c�W9q�$����)�ur�L���V�l���d���MŔ�B,��!��t��|Y��H\_:YUE�&�mu��x�J��٩��V��n�ď������(�ܺ�!;�v9�&hV�\�r�j�Ldd���C<��arȕj��ο�*/�ɿ��o���ô�--�Z��v�������2��>38��I~�W~��o)o�7���[�f����&X�<�����C?t���J����=~�W^}����?ftlB�>��x%�M_r�z&
��V
D)���:��->�<I��ܹw����o���d*����������ib���fthZ�ϕW�P���e�����~E׍g�<ý�,��,~_�f����Z�02�R�i%�i����/�+�3qqfvJyN��o^]#��2<>���P�^1[PCMl|,��#p��q�3�G-T�m���ߢZ*�r����´���Ɛ�j������N�z��Y�{�#~���88z^�ei2�T��>���ko��cj"D��Q!:f?����g��>��Տ�����|���8��wK
�z�6_��3lm|D�W�3���x�>C0Lj���k�ib���pom�Vo@1]܋����?J����t����j9O���G��������u��C�r%��VOP&�9���r��K����g0%��z�ln��O��l��B:���+W4=DtA6��-�>B!��,��N����ħY�ȳ��db�	j�y��U� ����L�"q����J���3<q��7V)�{{Vn�]�T�RmU��]��&�V�ڃY{L�cnX�ǁÏ��3���*�Fo��lYA	�)��f����Ĩ��X��x<�0s���y:���V�z���-���+X�������I��M`�KjG�f��h�VT�ͽT�I��Z�>29U�i��o)B�j�A0~�\3�����ڃd�b7@("ӮN�N��;����%`�(˵��1�����Xl.u�+m�uG����I��C�&K�/*+��֑!r.�~�q�KQ��k��XX�r�G�S���zH��?�E�Ż�yk��Z��w���}�{6�K����Z�?"��b�&y�1����1#�H�ZdsU��O>��k/}�H Hz=K6U����x�a�V'����94�a"&%����'��\|�/�u���v����:6�š[�/����.��D1�!��O�����r��U���P����4>���.��٢k����G�j�]�Q�^.252��fё�}e}]3}��+:^1]�*���d��@�4jv�@$1�:��{�.�n�\�!êŒ�W��7�}�Ό��M��4^�þY�pMV�b�.`?�{Qj�<�N�<��    IDAT�?��o�E�]��`5XYط�\!�N�j�������Y^[bz~RM$�kI>?^��6�K_�	�<}+�r�;�w���,�bx�Q�W"u(��x}>]m�f2D#])��[��2�tH�F�utK��*]����E�����)[��`qD�~�mA�]���i�|0�׭�dK����E����bQ:�9�)���4�S�P�~�+�^�x���q��y�:�F�t�y\�6��۴�;�.a�-��7�@ķ��f�w��*�<��ԏ�p�iw���dw����8��wX[z����4;n66��N�3��nӌ�h����ag ��)Fye���"ph�R���>ҊY���?����i
�}�g�y�����&�b�A9Lz�J�gx�8��O���ɝk��W�8y������u�_}	���@RA���f�Q�F�ӡղ�����E��Ztz?���l��W}��۩ٝ=�]	��Qjv���f3�'�h(���'���w������nD�K�5�|NJ��f�6:f������#��Qov��,^;�+��)�1��bk����7��YZ�K��I�S�Ԫ�u'�F��_�)n�x�����&�y������_����RnW����������1�<��w^�ܹ����u�|�=��F��6P$2zט"��0ut�.��&�89��`��^{_��@hq����/����566WUP��9~�Q\./�n����~�J���f2��-o�������9�� �}�ǋ��ebdJ-���yNj�:�G��N����ܥ,'O<�s�Q~PhH��tf�D4��o�I��c����D":�2�M�����r�оg	�p�ƛ,=����-��06�d6o����ٵFx�3���?��o�~��������㴻�߹I�_ef&�����&0��Wq|x�q����������[���t�ffO�ZJ.5�RHA3;�iIqhއӜ��2w��hw���W��˗U^Q��fN�#����%�!�1=c�Zm�� �]�&��S?��4�ο�"sq����$[ŢB�c6;����;����H��\�_|�v#��Rp��elv�B�E�oS>e�F3��Xgn8Ʊ�1*�
��Y�]�n=$Y����px\�pUC�]V��F!;��6�~�3��ռ1��)V�r��f_��TN����p�&���!ErC>,�*��ݱ8����^Z�ZO��(T�hQdE�Z�c��<1������}�q����ǟgs���U܆��]����V��x|��TJIqwG�łNrd�'Bs}'{-BK�o��D�&���������9Et�YN��ڰ�n���	�����drf��a/�����k���,�c�(5���Qi��\�v�-AV�9��3"l\�I��W�J���nuc�Vl��p5ҷ���������f�z���4�"�EYc:�j����-��0+k[L.�&r���
p��uVW�Y\Ͱ#�,�Ws�O�VM��W��|��(,�lcO�b���|t�6��6x��vk�շ� �$���j�P�q��m�8���8�.�O���l��n������~�r;�5"��0P7V	���U<vƞ�F�K��%]�p��g>B�����ō�W49�������6����>��f���"�p�[wohTZD�A�*gP�f�E�]"�[d:RTYmNm�^�%���BHV���S:U�4�z��|��*wo_�	����e��~�����d��%K�:��(R���S<N)�cjt�p8N&���q��a�W��2�h�j���W�B��Z��Ʊ�kk�r��Q����N��w�j�Ȧv���@l(�����+M���M�h�'FFqh�����*]�b���ť�,��zO9lVm���$N�K>�Qkl`]��դF�f�H�������J�SSSJw�jW|N��V�u:���x�M�#�z�̖$6��{��H�r���`] Զ����#uΜ9��?B�o����+��N��o�o�|a/���!݆LL�vU],�&���O��$���ǟ���'�I��?
� 7/~��cc|���K��$�������ςɍ�S"I���.|�@�G�<���]�`�1�bT�b�MKb*��Ʀ�����1��?����7_|����oU�V7��˫:�	������5ƃ	2y���4�v�i����o�.�QAz5����R��eԴ�F[2OWy��^,��;�^�������ݽ����jQ���fз�����3}�0�r�R>M�f�buP�Z�y'ev�	��i��LM:�"�PT#����!�Pjr���D�S��{���?��4j(��&�D�=�]�F\6+�n�dv�׌� /��S��4��s�U��~5v��{�7���*F��W�xE���}�����y<^+�=v�_|�?��?�L �2���[������C�Hm��dM^J�N�2'��,���%�'����o�گ`�[Yz�@$�������8p������􏿦�����|M;�'�|�ѡ/�_q��[؜Ufv�,�����A�}�%�d��Lb8�v:�n�(b<A������٠��V�.f:���J���q
�΁C!�mC��������c�g;[8�OLQs�s��c|����C�2���Jax�~�!�A�_������K���7�4��-�� ���OF	F�䳫=J�m�G�8=�ݺ�˙�����Ĺ�������w�5�<��ɑ�������:x��D�[���i*0?��.�3���_�g���ݿ�}�/^'UL��c��v��>͡����f7���
��_�����q���B%�H�^�Y��*�l����-v�z���!l�Q|c�fh��:4���bgkY�ʵF�J�F>S��A]�]n����e�Ǿ�)��e7Nb�$���.�O�^fim��D�X�S�U���v�߁��gal�}!��}Ӈ	EG�o%�(��ΰ�N�/F�j���X�Zā�j�X�f���VML8�<�����op�����KejC�D�C�Z�4.�UA���Ó��L�j�HL̳��Oq��t�γo�Iz{_�E�]�m6�ηXI�:�띘�1t�1A�Q�K`q�[%��E�a֯[�.��B�I�bfߏc;E&W�ν�%U�Zg7[`k7E����2�hf0�w�o���t�����I
��6x�;��jM�f��|���;�����2���Opzl��f8�ا�N>�:���#�|�����CǮE��-��NWk����*�"�n�'��7MlዔkV��_��d#��.�+�cC�9�\y�'�`z4L%�F}0��z��;D�զX�124��a��Mv�5s����,o���̑�(qO�ziE�(����#_d����.֮��
��vZ�*]Cc[� ����MI�����
����/\S�4��'��m6[�#��'4P���y��/���˕"wo�+�������~�^�����m�$tfJ�R��>�D�&�jE��5����Ĭ�>�ծs��0������j�h�4�$5�"�� �R�tr������c���S/n��}�������zt�"Ϭ�egrl�������������-Ɔ�����)��&{�:�Ϝ�X���'�HbDW�~,�!�n6��l�j��#�C���9|�(;;;�-�G�J�(����N��v���\r��rM'�"I�m�����1,N�Jb�]�no/1�o\c�cz�o|�O9r$D��gd����,�����?����e�/��gI���6ؘ8�84M$72�����un����}s<����6����4����>Tٟ�ٷx.��O}�LO����.�}�h��B���?���}��g�!����xd�\�B����c����ߣ����'?Ith�rU���,2;Y}��
�f�ݎ/0��y���0f�@��������?�V~+�Z�b�2���Kl�|�K?G��тf$� ���Y����S4J��}����T���A��d<�$_,����z�S�����Y�*~69�0�R��3�J��N�$�+�����7S���Z-䊻�n"n�\QW����M"�lx=���Hgr,on��Q�@,6�F2����}��ɓTu.���͇z����lUx�
��U��\�N�B7�Ӈ����.�����#��W�Z���9�/���M�Q�K�����<B(%�����".'<��c���G|���!
�(Y�9��eOo!-����Mb�Dd�Y�����>�BW��Z)�����5Fǆx�d��Me�aB�a��[���p��f����ԫ&l�ٝK�<� o���c����x��wi�w	��L$F��+����#Q�G'y�����?2A�c°����!z�	�M3���!�[k0�H5���ͳ�J�d��+�b4�a,���\��n���y:F��-��7�@�g��iV���L�3%��牎<B6_���_��v�C������pD�tX���[�x�N
���ٴ��8�����ٔ�Z}�b����ǧ�_W/�qX����m��+s����s������>����u�� �k��[1[T������fkG�}$R����<���%�%��#��#͍hzC�f�b1���KK��!*�<{��'���S�2Ը~��j���7I%�h5����x�a	�F�b$&F�X,����}|�G~�c��?���_�+6�0[z�+9�F3�bY�J�����͏�����t���b�8��׹x��-�#��*��]���^��t��x��D�kgP���1���<��>�N�ȟ�Y[9���03�j0�Q�x�	y	���z�G���7<�έil��PO�u;0�{thh�u��`)]� n�f������t,@O�>��j����` ����Gc=E c�k�`�������ɵ�|�[���իD!���_�>�k.kg�����6�1��\z��<rhO|�yڙ<�k��a����>_���N���n0;��i��M=�lkQs�-���#��_�����	���[m,"f�5p���3P���,Pb�ś�6�� W��S?K�hb���t�;*�=�nj�h��eM�ڧ^�e��/�pmy���IM�H�oa�wԥ�X])p����1�x��w�c;2a饘�#�g��/S�N���:�~:5���:j�}p��'N�|���&筛�x�~�\5D�4�Ri�/��/�aM��5��$�ii���#�j�I�w4Bt���QmwbtD�EG.�?&F�TS(K��T��<:1��X�"�i7@/[�T*E(������,i�pO��m�~�M��2�s�$w�H�l+�(����eflLs��ݾ��̴j7�9Y�m�2�T��M|��G�"a�<|���f�4���z�A��SL�DCJ
����m��V+�zȗr�"!m܂^��3d2{v8p�t&�7��M��8Ɂ�C\�p���vx��>�p��?��Q���NOr��U�;��T�Or�ʖK������C#	ݞH�(�ȷoS(�����y݂m�/�T%��n��{���gOQ�4��EO�Qsf���ݷ�k�����X_c$���_���r��#g�������{jNiֳ"��op��q5v>��*�z��;ݼ����?���a�~�Q�|~;��Q+�;j���m~��~����g�p��I�޾H(b��o�������a��1�5��ސ�Ӳ�MO͓ϕԍ-w�|.6��;��/���?g0������O��k�w;͇�}�SP̉��j�$��&<tp/�i�D��� S�E��'�� ������!n����d��vb�Ke�^.����SG}���7�\!��Y�q2�jX�q\kpe�d��;���Q�K�M�Z�DX�[Tj&�&(�VX[�ҢP&g����`�KWn������jQ�z���l��9�	�F��p��-n^;�N2)Z��@P-���CaM���O=���l3p��k����Ϝ=4B84�s_�-��[o���.�M��Mk.��j����Gy����%E4�&�$0\�0��������R�X\�,�!)��E��&Y[���r��f~���E� /���]�L��!�M`��ؿ��wA/��'�p���V��jW)V���I��qLO����t���4
U�.�*T��>�B��.���F��5Ѭ8��/p�����?�.���M����a�"ڴFG��?�� ���S��׮)�3'x�?����z�?������!��fGǸ�x�F+��ѣ\���#O~k�Ih��M�����^=Ð�ʺ��"6�/��)Qj��ņ���W�LF��M'5��l����,޼����Vk��.�f�K��cx�4_�;����bq`귨��@��W���!��k�	��f��G�.&�1��2�j����N#�\��G�Ô��6��H�e���|�ͥ[�L^�=+��=��~wȣRK����xp�-̃2f<X���؈�q�m>���&F�N1�pD����+���UJ���/�ˬ�ϥ�Y�X6����Sz�Y9��0�ó�f��=N�ޡ\�����"Kn�6hck]�B�N��B(�\��ř��g��#��Ln�f�jw��}��囪�o�Љ�M�W��m������LL�O��20=���I-�M��S,��p�����:�X������]}7˅-��'�	�-DL.m^��m ɋcpЧ*X������T;^��O�8�	�v����}rkK����'�'>:����m���
c	Qg���;���K�ѣ��1>:��ps�.=����~:v._x�j�!��fu�:��7���*�F�8q��r��B�k"vQ�e�u[D�15�b0�dIb��-,�F��)0�䣿@����&�v�jA�N����±�6vG���@�8�:��,&��f&�~������
��r��<������ަ��h�5�8��5�k��z�ݥ��%��L����/�l��|жbn�0�B$0��g�y����l�(,~u-�+e��,�nc��7#	Z~��^ήϧ�Č�	e�����$�I�Yi e�'�>�~�G��ҰKsn��� (�.����"H�sѾ�R�\*24�R*�,J�[�Y�!@��׋_��7o��n�T�2C�0c��BJ73�r���H&�������<����Xcl|�ۣi�������m��7�[����,Đ|!����PB)G��i���SS{�nK��?|���zJ��۷���Aaa���ӑ\l	20���ޒ�;����Q�2Ŕ�M&����"4�02>�:D�F�-{�^���N�v;p�-l�<���\��"��?V���ccx4�'�%12K�ץ5����*7.�hn����v���?G ��.���g�}�o�q�-�w�L;��
_��O�o��{��!V�6T������:�\����9�'��fr��}�z낞�W�]�\�s���gI$Ϯ|�.ޤVnq�3�(:b��F���h���tp9�ڄ	״+�}b�|�����?o0�J��_���xR���_��R���H������f>M)U�'R����}vwRD�q�V�X�w���N��V��iY�jS:�V�N$���o�;9ud� !b����$H�S<��J���)7�<]M�X,���s��v�hT��ޭr���i�}�����Mas8��L�.i�nt�ZZlAf��b��㘭>�(H�e���ըc�B�Q�T�x,��*�rCkO J���;2L�$��
/~�0wDl-��'���c� k7���$k�<k�<��1�_~��V�d&R�=(���0�N�jt*�MV�6�Y���N]M���w��q�=
�3�ڠ۫��-
ie���Qʅ6�#3��^Z�N}�6K���?8A���������ߦo��ؓ_��ӟ�w��a�fg�&�R��{˴Fz}яH|�L��<��c|t�C&�|��_��������
o���n3K���m��"#I�`�u���|&�����G�׿�G��6}�^z�_Я-�ȁa��Uu�ˡ���X^_���=I`�y�1�)�ݡU^�^^�UI�V^�2c�y�?��F�G�c����    IDATV�+�_O0�$�Օ�ْ�1����{\��U��_cn4�BapWh�'?��{���j��j�]b�ҤK똜����4	:�}r[�
A�Ƣ4�5,V���jw�g��{�cFe�ժm�vVŇ����ɝ�����q�����N�j��$�XjE�/��y��J�liG'�_�aO�o����Ï���D�5P�p9�]�X����Cv3�8�v�Tm�ԕ)kN�������ng�VMP���.s�;�/hn��6o�l!����D�N���c��܏���0(%r�O.�ԢA/$�Ut�4@nW@/�f����dz� ��<F�k���&f)RٺJ~��hs�ass����`P��;��4ӼX�򻈻=���Z��5�f�� �A��tJ�L"杁�b�M`�g���`#�䥗^"h6�s?:�����_��2���kN���cl8h���u��+eފ�0�Oh���;���Q<NY'f��w�#�O�s��^�6��+z��vrLM���Y���Gvg�̈́�� _,�,F�Y\�&M(�k�&p^�sp?������m�ͯc��޼G,�bks]�[H�hn�J-3��R���Woa��0�,loo079Af{�� �Oe�006<�������q�c�9��D�h��X�Ô�)
�k�u���¦�}b�Y�&�&���;�gx���x��+�L,��D)V�8�(����g595C�T����
��Bٲ� B
d�^��R&�r��VfldDM$�YD֦=ɶ6Y��1����h�(p|i��V�N���Ϥ����ew�M�K�lZ��������_W�^��ts��U��0:���x��!��E#uI/���/�Yz��T؃�"2�0�qy����B&��d��e���'�=덊�%R�&�;�7�"�֭[BA�H��H�4�i7��;Q��r���ܹsj�Ko���H�r��g���$���Eox��eb��~�~��ZC���3i�(ZV���)�zrΜyLMh���h7*�-��I�"�x����1��駟�l�����l뱽�KyG<	6$����=,&3�?s��#�tb~�k�n����Ѷp��-<>^����!��������fg�����a�]�������:m��^"_hOr��U��_���>u���K�J����ꎦ��Lh�B���#z��>-�%�utd�tfWk���������o�����/��������)�^�m��E�V���`0xp���9ΩG�SW� p��6i5��Y�+��U,�;��Qw(V�i�\�b�R��q�ȱZ�<A�S�u,I�g1�����/VB)�R����b2i�z��������2DQv��4D�,I:݁B@E;#j(�j�ht�C ϝ��uL/=��ct�rXv�<�l�ʚ� �!q#I� )\v%Zc395�P��h�Bm�ZG
�^�qa.�.r�D��k"Cl|�R]����m��+�||}����b$�ivc6�t�i�#m��N`J��4��43;K�YӢQA�#ͥ�ճ�w���v�r��eU+����UۊR�������e߾Y07��>�u�H4�+8����Dc�4����̥_�m���$��U3l�s���<f]��BC�Fg@�D�b�b>��Ub����akc�ݡkc��Ja�Y26cbj��铌$&���6n���nse2�L�g(dEo��8î��cL�z�Jǫ�q��C��bs�&�z���q��IL�T�\R�����nvj*i!��,�1�֫Uj���������o������{�\z�/�R!������h�O*��I��9x�\N��
���RU`�F<��t����ѥ�N)���S-�p�z4�-�ȸC,oeH���z�F���cn60 9�º��g'&�\�r	����qY��N��ԥ��ɑ8��:E��K�dڃ]��DbK�2����(�ڪ�VZ�x0��d*���Ӹ+�Q�U�*6�&�^����Მ�9��Xmh�``ܒ(P-+�KVc�JS/)$噓	��#�m-��wX��[}ܖQOGY�a�DNU�\��uY��XYͫFkv� �v����m�w��f�����������r��7��*X�.E�4u*� c'���1J������tKy�<���S����&y���?����0�w�Y)�$L�E%��O(!W�k2�#a��)�J�B>�\M�f&��*<��}:�չ�?p�r�̵k���T��6������B��b8�^֣�Ág�4��̠��Щ��^�h���v���(�HT��
�����`�6)ջ��nssi�@ة��l�Z�cC>|>��ԅ�f����{r�^n[qd����O��M&�Lj���$��d�W4Db���|��%D��������mVW�t>�m��O����+��o�bQ��֨[VV��ͭ]�@���Z(��ZDȄM �:��ɠI�0�sԊ��ns��K
�z���12}�er��!��Wke]Q�W��Lv��顀�%�T�qw�~66�U*p������*�iV��&q�l�*K��\�x�LV��vg�׎�hbww�թ�vY;�\:}�I���*��	��N�g�X\_Y%�*X_W���w�-ؑLh����%<�߻|�?��/�cw7�zĲ$��.��tiV�ȡ�����sݤ<�����"�(f���P�N}O�+{rk�cGg�x���u,3�n=�is�nssk�}�'	��d���8ƁS�F6S���-\~/�`��Nh4�Y"�]�V7��\�ޅr��N�� Sc\����8�|��Q>��6�\�����e+���ms��"����Ar�[��MF�b<��c���g��9ZZ\�aN$:�I�u�o�G:����U/��c��lmmk�au��L�����د���ZQ����?����W�7��zOe�v��51=}����_������{���d3�?���֦F�f�^K4yf��Z��M��bd�.�,��A�'챎NTt:�+��i���barl�)7��:O�$I��S�h'�UP��.msh$�@Q�vj�z�f������cv-�(�Z�#�4�e�&�F���Z�-=�p0��l��["�	b7Ks�z��3b�ݫ��Z`�ɂ�ť.w�7B�lb'�R<�~[���E
u'[;E�It��o�l��L&�r���N&i�&�rL���m��4���R��y%�^�F���7b6���0��oi'��Խ,����b�P�l�qu��Iq��s|�K�D����qQ.�U\%W�Yi�$T�%Bj�߉��VdH02Gfw�ZMxU���X�f�b&I�R���20�t)_��z�>� �q�B�,~�
[zmz�M��N���P�N�Z�ߴ�����4�
66�blT4L~LV��v:�Eq�����^lXg`�e�13:̠ՠ���GU��8q�L�`��t��$���l��@G}-4��iw��F�F[�o��Ѡ�J!��nW�L6���l��A�.��,�X@��&;6��n��}��5�
$Y���璯Rb�8d���^�r�����g�V�I�e���8����>{�kop��EN�0<���kw�T:vKULRlZ<��}�w;M�uJǲ��?j�[5˵�,��Art@ە^�0D}{Soc�^��Z�n�H06J*�S,F�עߩ��r���9��I�c�z�KIo�jO�*f\փU~_�"?���p�*UbA7nG������d���X�t=޻q�fǀ��Y��1�~;�n��+���db��p�z)��g�b�_7��o��(�JD�������k�1�9³O���x��W�K�ij�����N̨!S��v#��͋�\�ou���@�q}a�?�:)E�����}�I̘�:�b2�Y���V\cP[�ei`����#���Z[af8�H�G��C��W��h��/+Q�zʤ[�'6��j��}D~gt�����u�C£a�g���$�҉��&����Xbf<��N�L��N��?>,41�[�NM�Y��*�Sc4*��]q�TkyN?rL'1/}�E��a��'84Gn���w�76p����bH*a$�&��!Sy��mC�7LjC�4�E�_8M�1�G~�gh4�X]!��H���뭒ޗ����?ĥ�@��E�n��=iv����f�:��D���Q��u�"��|��t�-0jm=MfZͦF��;����Y��F
�4.�����w~z����gЯS�����e�����}663$7�ڴ<4��i"�h����&)	�rtT�{Z*M�sj�ݠR,�ٮ�J��<+ć���$SI�'�uB(��\.�s�=�r�<:t�7_C5���V�^�:��(��+-[�hTנ�b��l�7n\���r��Q=�d��$����!r�����@'��.�`nfN�K�>��i�^�"ږW7HH��١1rR?�Z��u��k`�Um��M�J�=6�s�%���.�����Ń�ᬔsܼ�Hll����|G?�GY vZ�M�I��lo������D���7�g{��"������˷uz+�}�BQQWRV��~��@r�%�H��q�<-V��=�������������o�>~���Z�p럈7�Y�tR��(W�df��1��?8=��q��+�/,�IWU�����L&�>rȷ�e�A7C1?~�8�*�g+�9R�ɛ!)>/j>PA���7K���J���؁�jA�<$��tDf2�=�Q��K[Ň�8��F��')%AR �����ez(�C���u��(@Q��WK5u�|.�f7��լֈ��:�
~|8�N~G��"�}���d�MS�7t��d���w�� A_�r������\�&J��j��/fs�nG&%{a뽎��-�{��F��Dt�ը/HUV.��e%����\�� ,4[#66��I�[�i���*噞�\���g)S���|��/s��e�:{_��F�3B�ӣ٪I���!�=n��pG��M��M��g�3�kդ���`�a�ۨ����� �65IL=n��F�L�&�Z�t:� Ř#.6�Ӭ�l���C��H�����5v+]]��-�F�E���p=C2��B#�spr��ˢ�S���K�+6HnW����ڷ0��%�u���4�@��fI_\чH���yt[��y���8�l$�\����n�ȑy�Q�ꅆ1e5���8��&�l]A��]�O�����j�FZE��� #�lf�,���f��#�!�x[����fg{�g���VV��L�]}F���m�>�7D�?P���E�p�FE�㮰�&\Ni&:��m���N�t��5�VMxZr�v$;]P&I�b���}[Kf�!MW8�,�z��r�U�m0��ؔ�L.��Z}ZM���&��8�e�)\P�]�qFz�:N��d[a�1�H4���mX�VRI6*5Ʀ0���@�sd��N�VPⅹ�c����FWVz�u+wW)4�D�&���v	;�,��"6{����?U����W�>ė���3���/hDY��f{�&:xf:&i���nѕt��l���gS#�H0�J��Amwg�ۤ[�^kw�d�3ƪg���*V�ѵYK����D*{_}~�*o@�L�L����I|ǾW���p[���Ar]�w�N`jd�~�N�����V#��z�L32=C��W,�H`d�P)Ʉʌ�favvZ�?����l	ىE��euiQ���gImnPI_�fHc����fYeRpՊU|V}���q@�c�eec�J�n�����y�O�L�A�JP,V�Y=�����=�p�ʥ�Njj������ڈHȂ輽��p� C�X��k7F��a��C���,�|�wA�dB��{H~�K'b���!��]��Z���f���wS�����M������E^}�m� �nG�N���c|t�յ�_��C�` �frK�8i����e3#?߿��ߋ �B�`(��vR|
Cֿ�2"�fY�J�'߯�odc���Ĺ'���"><L�R�5�|�W�\a$1�߷4�2Q�fZY��2�[;[����X$�����nn&��g��"����˷�Me�T2:��Y�U9ۧg��`uS7ab�^ch4��Fyn�GG���h$��K��crv��en-n��Y���c<����׹~�.ё9�+/��	ޣ���J�4Jry9I�)nn�|��ģ��$t���N>+zR��[["�p��'4e��8��u��Ln¥WN�����+R�'����;?�S����)|�����j���,=z�X��z]�zU�V*��n�u�\����K��+����h�m�1�VR��g�n3259�Y�:�6��< �6&�d B�.���I˪�g�����X�%*.�~���$�R�@V�m��i��IЌb<�^ٌd[����nI.�d��n4j�hs�5��ڨSoI�F sߡ�?�#Q�R6{55�H��q�)�K�R��V�R��(Ѡ�*����f�
��6�j]���C������0Jq���t) &�fhԳJ��չLh�MAa���u�!H��*��,���0��S+� N$��'Or��kl$�R,��v[qXt��ވ�*���c}.'�dG�ȣ�N��ڼ���ߗ)�Y���y�u�bi�����l����%�����ͣ�R�&��������A��w���̗�}וuv}�[wK�$˒�a��A��g����L0���D,3��0���:�c��`c|ɶ,ɒl-u�������ʬ��/_��/�Ϸ��M�D�"aK�ՙ/���>���s��R��!� ��9�r��"�f�#��=�0�~�v���DR�d���-lo����eW/aa)���6pX����h�p��9��͉V��nA4�%Wqan��Ԋ���d�n����%a�8��x�,������I�)��Ò%��ؘ��A�ב�C<���,KE�������	�v_ �#��6�:�L ϡ֨��*H��\�}˄7��q�Qi�`}Fw)���ehZc]��;<H�=��v
v�#�z� �wK�{�KG�k���+�P�6a�>��M[p{|һ�X̡.ݦd8"b ��Vjl���+
�&5�n��X��6 �X$ Q�Ƣ��㏉�h@�|�/l�t~������D֘���V���f	�o$yg>wH��CWm�~�6Jx��>��(����4�V���4NM�b��-13$�~T�>J���b� �)��A����=B�h��ۨt;⮝�g���1-�d.|��ß��KO�lf��2籸|�F����uy2�F.��z�:B��T{2���K �����y	�VG.�m�p�=�����n�ho�K(�J�VK����ȡ���tċt�����ѓ� ��_�^��[�Ƀ�@Ϋ�?u�1TQ���$,8�0
]Gmy��'�5 ��w�x�S��cD'�ǋv[��=���DI: �{�ޒ���[x��_G@30?�cVa����p��Ǡ�;h���� pZp�,8������VG�/Eˣ�v��R�V���
Z���� �pٙӸ~{�YQQ���APx�=�����H��2���:1G�@tѸ�\V]�j�D7O���B�D���PD������0q<Tѐ��|W�z�άᑇ����2������,��s�M�Q(�Iv�܃����l����4���#Op�ڻx��נ��0C�=�xH$\�V�h\L5���gtla�
�C�/��7���Q.U�����;{{���Ň?����/�Ν;{���#	\���=p߃x�ڻȤ������$˕g�j�*C�]����ɆY�_8�ק	y�E�L�Pkt�ыں��[��g��F�2���>�tw7�$n-�I��>�Az�D3�{X�k��	�sR�Yl��vP�#Q�&��ӆ�Ա������T����}��8(UDW������޶L��-,�݃�����L�b��~
ְ���=�V����^������ucm&�$Uǅ��m�,����j��@4��⡔1��=X;.��<��!f�q����O�������}���?������K�W�Z���ۍvπ��qx�C�������s�v��!6��B&z9�u�l�`��T$�TD�CIv��'���7~2#yؙ7F����HD46V��ǋ�m-    IDAT�"�i�V�'BU��P $�z���թ4˘�O�bԪ�Ee|
xP)������ 	<�O�^1Ǐ�3�P�a,��)�̪U��^�,�w�0q�-=�tB�ъ�4#��:�1$��+X"z\���8��Y|�ٟ���e\}g[w�d3�(��<F�]�i6a&4�p�VT��%6�[:�M�na��A�/���:�c�Ξ;�௿�ad���$X;͢tx,�J�^�l��!��d�O<��ａ�lJ�=�x���YEIjN���Y��Fw��;�M�q�f�i$CA��3O�����0Fd��a�D����P����>�L&
�u�E��w�ˌ'��S`x��e���vE�|��Y�
�o�Q����4&	qﾷW�^��\fW�1��q�/�	��z���nl��hQ��&sA�=E"� �K��`=X�@¡y��-~��<ı·��_�6����q��#���0�{hn�� ����`�1Ǡ��Ɇc�`t�L�T�>P�����{֤�bd����E���Q�D#����F��qQ���h�/��1B~q	��>�n��w���R��P"�Fǀ1"���bqv+kn��	Ɔ����|��e��жa[4|i�Uc�t�b,������O�'��*� ���F�X��ˍ����l�V	�4U���#�{1��^�$s�a~�Ze�F?ՑS;�	��Ʃ���U"�V����z��ipJ�&��S,`��Pڔ��	�;�LqV*B������r+X���k98�S��)vj�������&S�2vib?�4���vzc�V��	{Ї�bޞ~�&�����]x�x�	dfO�+1��,����� ���F����%P��d�!3��(�o`m~a?ߦ n�3��l��12]��^2d@<�<�W��ץ�,5��j�����<�4����Ĥ��j"�Iw�� /�Y�L*��ㄮ^Ց�LI��I�=Bq�6޻
︃|��҄{\E Gr��#�_�e�Bq��ә�_LŠ��K<=�i �>�f%��^���icfa3��}T����AE*�R�1rp������ꊰ�t�rb�v�̓�* �׈nw^3�̾�/d����CG��	S61�z��|~ZX:.c�v�v��Mw�[o~OdQ�?���x��/`��v]�d:&T����.f	���6�}3���+@�ΝM@�D���#�X��nm!71)դ~_���R�ɞ@��!|�'y�.a�*��ZY��AQ4l��>L��U�p$�C��\.y^9�er4���8���I�G�dH9A����u<��I�8��3��'��a���@f�,`w����X�&����Y�`���ј�hO>�!������j�&ʇME�X��ұ�{��ʹEh��q�!QC�}��*��ҋ��~ݡ���Yxl
;�#A�*Ї*��$Å�B�D=tz����n���N�'�
�4$i�l�p�^��#�ʹ���Y������v��lw$���t,��f�/�;1���}PU��������/��oZQ�����o~�ӭʻ�Z�V��H$+.]ǥ�? xscg��jY����O���r�`�x���	4*��U��U����1�Q�q2k|���n�����'"ԁ)BX�Dd �a�T������s���wXc��ƺt�z�q��a�nS��Q9�@"E&=�.5R*5�r\� ����ԒH�OJ�M���x,��I}�vۄ/C��KU�Q��I�4��E�@F�)�N_G*ˢv���0uC���YC)K��bp� z5t8�1ج �����QQ��A�c��l��m�q�[��L悧T���<0����H��;��d~F�>��&&�E�Ǜ��=��}���!����"]P��0<L�(cDC^\^�A.��mCC��t:=Y�Ȗ	GQ�*��;�6^��#����\>��؆�������2�Q`��4� � �o�-
94�� ���￞��]���ug��ǘ����o!����7�q�J�������H�C��Z�]�Jeپ��4��O�A���a�0�4�
�m?�JP�u|�'}P�Mx�����������k�[���vK� �W������>��+܂?@8��]�@��Yp$����Ebn����q�٧���1��b���H3���g��Pi긹�D��5�4��.�X�;%�lө��d�bluPk�o�5٘���[�!��'=T�%�0f� �x-"�vJ9��Ɗ�*曒�+7o����x����;[,�atMq�S[����[�S�(n��HN�4����Ú����Y¼x��S':���=�=F~.�;���sci�!��@?��B�N!�KB18z�^�92�[o��l	�ͥ��M�04�0����j� :���X��v�%�\ݎ"w�9���S�7��02�����J����Wd_>�C@�Qݿ�Sɨ��C��2�d}'�a:�z�Q�:5�R� �L�ze�&�-�j��w����]�i�M�� q��D�ˠ���&�y�Rk]�[hcx���ч��1}�Y����+`4T�|������!}�i��)<,a4��n4�
������{H'�'�7��Zm~o�X�0�h���ZHGX�	��ڄ�@n�I����W�VJ��XdGf�Q0}~�]��:�y��z�F��Ar2��SgpXjA��έmh�8�Ju�A�>{�.]BZ�'k�?���i���[��z�2�����'�!��u�3�14�%Dԓ 2qb2+&%n�����_�ꗱ�4�������qjy�����8u�<TD$�������$�f�D~W �{{�!��S��őH��nבI�d�J��,(�N"�����4�h����ף�""A��ClM�$��QO��B��d�	�%N��VS>#a���b���!����L*� KՊ��2MH�����"����'��q�Y]�_�՟��em�H���utڜ�D�H	��L2#���t2�o�F�7�ell� �LE19��x��T4�[�oa��_$$y�|v��8{��YY���z]�G����SR~����3g��T����z�/`�?��ᕬm0�=��C"�r�2�v����S8.�$읞������Ti��9��:�����?�;��_���(tK����5��}�~�[�4�/�O'r猒�h�T�a��(��H%H��E�yx�����^��.zA:޲�����,��Nt���4����^P/v#��|j��$�������ǖ j����C��C A�D�D�^�j�0;�$����8G�47t݄[� ��G�����hv��52Z�C�c� ��Ѱ��6�����x4p6$��)��������
:4A4Z��`?��j�E�7�Nׁޗ�?蝾|��B�*k� �Ӥ��đI4�����濠�#��@�E2��Jml�|��AvW��=]o����߮6����﷐H���+Hl��.�^
���	�E܆?�ۛL����m׶$|���ʅs��4�����Tz���#e�>�>˖�w�W4���(�f��-�ԋ�*�E�#��P�S�m�yRh4�h4�P}@"���j�҉�U�cko�t
����
�n�G��Ǐ�Tg�a��Pi��w�^0���>��T�T��y�~�у�tïy��#�R���>�1���jF�g��^���q�D^��ɤ�q��Z���S�����Aш�S-$ݜ�-z@�6G��(��ޮ�ȉ\v��C����N�5cp܊%cf�ep��󙡺��~�m\��=�3Qi�G�����.���p��?l��Ɇ>ޛ~_H\�<����T�<`)���dw�n
�����8��z=�c�zK�<S�����H��,� �h��ר���>cM�ej���D��� �!Lw��ܧ�t��ѻJ��/���ۡ[&�ݎ��8�iAL&g����y؊�28�T�DeCu�M8F����?�����?����_D8����0��0���{6���~�Y�$�}�>t�X<n1<�y��c�������HCD1���ƭ��z,�L �v���U�"�CX\�#I}Z��SG,0@�p�jM�Z�!�a#���t�S/nB7F�G�XXArf�U��.4-�Pb�6�҆�d��4���l��w�miR.��+H����)�P(6'�wXq�;-4*;(��H?�L҃l�Y��
`�ԇO�����o�o7���1��'c5��%���E�V�&�q��,����1@fjs+Ĺ�_l�����#��\]=�ӧO�N�@z~aV؅B�Kr?q�'#��� 2c2��	ɇ�ǑJ�ed����ڙ����z���/�ѩ�	��96-�p\<�����A/�Q/���ߏ�����a@֐�7��N��>|��	���8ң)��׿�tfRj9i"I�ߋ��́-.��<�|v	�����!�)�iao�Pܾ;[{Rݗ�Nb{o_��b~F�\�	n��XC F���?#��f�d
z��V�)`>㌼!�d,�E���F�[IǳG�J�F�]���e(�)ϯ�� ?�����pi|>8����ܺ�|>�lzB����(������^S*BY�ǿ/�M`l�pn~�b�o� ��!39�_}SsI�y�U\��ħ�0@Cd��hX�?��K��2�N��R��P��,�:�	9���@6����c��L8O��P�"��J��=��슌M7,<A�!h6	:��Ѕ���ȿ~�S��7�o5w���?߮���A��G��6.<�.cC��Z�͝D��C���\nZ�O��%c�x4$yp_�#C��p��PS^0��p���P��PY��.��.έb*��.���fwv�$C�����ao�x�1�.l�x��f03�E�P��y�����F����*~.�G�+~����u���M�q�����:F�`�(���t{ZC�%��z�(5 ��1��%	�=����hǪ}��E7��$,�v��h�1��1]b��q!ɰ���`�@q�BF��QD�ʠM�}}��ՁT��}Cn�@(
��-Nc60<�J�R,�{��GS�0�-�6gln"�ߐ"t�O#��`=� �AG����N����c���)��'��2���3��]8�#��BJ���.O�ԙ�6OF�~��춇�I	�:T��D�o����b����Fh���+q�#nW`b$#�T$��k�P����:�^B8�|
I��������#��^x}Q�]�����ƍ���,�7��c�I�J�/�Y��y�m���X8�dzV ���.&�~��E��H]2i�zlJ S�	a싣I��E�R�G0���d{z&�p*��T�2���c�����+�~7:��H�l�tO������02_gn�Ӆ��<�(�<���@�x�cbs ������_�����Y ��n��A�� cF{0R�/�7O�t�DS�h5u��.>
:��ȹT2Z>a_h���uF'=�t7ss�a�,GL��#U�St��]8��⸰�d��6�<.�����h���m��z�!l�F�]E6�|v����O!,��(=��Թ����{�/�%,?�,���M����m�u��x����q�tJ��Jѭ�a1�P˭H��^����
�ǃB�nJ �N�D6�@�^�y .��W��'�����ETk�8{���\��:2I�nU���Ĉ���Z�@�>��P�D]��C8���S�����ݫa�4����hȥ&���FjfQ�yñ���F�x�h��D���tѷ�QE�|2=%`���Ъ��:�֭�J��t��#�p`�V�}UA��W��
��ҢPF�Oc�qMF��X�� ��e�U��:�K��>Bfz	�/?�won��2���r{�(A@C�M �x\�&~\W	x�;ŵ�k5�����+�}���PK&����;b@c{�t��/H��%#�h����x��z�����D��n\�\Z.���\M�M��<t�e�
�pq?��x饗$�.5�ŵ��\�祒Y�w�9��#��=����x��G4�CѢ��ؖu����N�O��z��j�;L���$e{~�1$ %�42M�ZZ���?�}����w7�-����ni��y�H���ŉ]T�FK�I,�e���
�43������{ ��kEu���L��'�7�n]�+�d��G����iU�����XH�p������I%�2��۹�e�4E뛟�Avf
���=�>�ǈǸ���\�|�y�-)c`0�'�d�	y�ຼ����77��~+�gF�ddQ�J�����MeAoH&���1�O�#�H��'��������QFa��������ح_��`h���G!��k<������gp�_��y�lt1��D�\C����9g�>��P���P4"7:�c)��}��"�p|tr��w�D������]�
�^���\:�����sU�N;} �kkp�UCC�9��K�O]�`XD��$rO�K�a !�AM]�{%ˏ�c�{?G��D������' whs�>����1�/R��a2�IټȨ��Q�*U�MR�S���t�XC	�"�ԹY0��'�vC�����!�#n��[�6E�<�� �����6r�ݣ#l2�yX�&�������uZ5�S� ���x��Y$�vo�c*7�1L���TI��8�:=q�i�J��m�c�ށF����?�8b^N��\�q6U�4�<Y�{$���S9M�,*#`ld�n'�v��uj���a�nD�u\F_�Vސ��W�^��y�o���{��R��<��d6�J��ۇ4z'ݶ�pWΝ�:�c�#�_���ES��#�u���UݰMƣxEO�qt�ah2��A����i��7t�{��υ�ރ'�`D�"�dm�ȡ1B�*�6����i���Ca��ȟ~^�±Ы���*�����,d N��/������GT��&��c9���*���qT� 쳡�R÷w��`$-��81`ײY]�E\��ýn_�w
Х��!���'�E��B0�R�]��:�OM��TlåQC槉�,����0�>�W���^��b�Ϩd�\9Pt{��c�^���Hg>M�VǐMZ����V� t��<�>�ͣ��ǈ���@*ƹ3p���@���X��9`[��C8<�,�f/��
rgqz�<������W����GG�?Kp�t��l����yx��0��[s�2���?�Y��i���)���E�j���<>���y�|�����M"q��sr*/,�;o���	�2������	b�x�3aU��;8h��19��j��R�]����AI�a�/]��v-�G�x�; ��Q+TqT$C!�fW��(١��b� kIMX�kg/��Ua�5��@���nu�"Y�;�b?����G��U�.������uq���~����@_�ĝ�-��W�蚈�'pks�'��>��d�V�1�1��'T^?u��  �zw���%���ɧ��2�d��&&�tE�:��Sˈ�¸���n����e�2~���{��7��t&) so�.��6굲G���q��1� Y1@�5D4����fg�+��V~�	9\�s�Mqc�^�5~Kk+X�sG�}|���E���M��ׄ4�(��in�3�:�a�B}��o�<�p!����X ��l�ݸ&{#z:ݮL���{:!���Z���qtt ����k ��V�-$��A*�*M�|�x�J����d���(Z�lm����,j�������0�R�;Y^\�շބOV�Oc��>̑
��P.��h���A��U<~������$SrX��pL�Lg斱���$�<��	��6M'��K`v:�A�Œ4YwvѢ\��C��o�)���r�d���w4�S9��/��{�R!H}=�^��ga��'��P�A:���x����/���ht��?�����y�������ns؅��1��2�;d�K    IDAT1'ol)�_�C=�
M�>�ر,ڠ��:qŲ��`���v��w�T*ǲ%�*�C�t�K�1��A��)���tPl�Q�0��e�S�;�]�j>���x���&�Pnu��qtx(����$��'=�ñOc^��P}A?t�'z�P�'e�.�m�*\̲c^��<�')�#ژq>�U��� q0p�ącDI�ח�����h����&`��R5�[�z �������5�ǚ�E�I�6�%���8c�$��[F6;���ݬ���߫cy!���D�1�X���q�P
���&k�q�df��L�j	�����2�q���L
�bI܎�lF�^�IW���㑀Z_p��n�U�qPF׶����ҹUD�.�=��,�o1r\�0L�b�^�P7"af��E{��hMǭ��1`��E%��t�*L����A���D�gB�`� "rݴ�uP@�qB^�vk��Iq{<����B��{�J����EX�:<�el!5Vd�U74776��aYTW �EC�*|T��@p]#v_/)�~R�k��M�-�4���1.��+�0����5��P���x�9t��3�q����8�o��%XF*���J+
Ǔ�h��1�QF�)�f5�/`�� �|�g*}Ú׏��584;t�U�*Z�rSKҪ"&�A������xٌ
	#H��L��8��v�F2҆���%,�O�!����a�rK�|qo��$B�	��ٓ��Xׯ��[��	 �!�̋I�P��lʘ����^\\�իo��g����4�����z�����Hff���Pݓ�G�}��0{5����	�a��w�yk���h�Jr0]ʝ��|G��4��F��s�����e��1���G�p�}��Ww��/�9��>L���߾�p|�*�s1$7��C�(���9@�*�y<��=:1X�G6��p
1O+sӘ�`:�]:��#�K�nSq'q��}����&�^F�X0{d����fKO�<��r��A�z@��j���0`yj�p76��1�S��k ����O���K���CX̕ӂpL��p}����p�iIQ �V�pKK+r �\ܽ��a��M��cdc���ɺ��~Ij�J��۸	O\�3��X���
�c�thA?���Nϋz=��}���{����R�Y(������̒hy���i��b���0ٛ�_{W�P4yd�hh�nc� ���)h7n�Z?1�y<��C	G�{Ei�`V!� ���忓�g6�~O����iT���n�I��1�x���dP�3�ͅሇL~7�z��je|.9�����{��ƗKg�J���D<��Ͽ�op\)#:==�A�D���֭;R���A2�=^������sнNH����MydS���$$�2)��-���>Zo5�87/Q5,k��#�=I�G��"S��Me���6+�d�8,��@7-�f;O$D��������Apfr��6چ����ⱐ�LZ@!��~��+(����<����j#u$�b&�D:�a�`Z*��#����O���Y=F���ӫ���H.���s�g��^~�e,�Ϟ�&n�r*Kaf~�n�F�ф����_�{�9����R����?�3��?���������;@�?��n���x�}�0[�N��d������D[ ���@8,�#1<21��ez5z]R����ӽ'����
���^)baj��<lÒ�FFDP�?��e�6��yh�(�	�K�kh�޳ga���-�w�0O,ǘ�H�fm[tuRGD���c��M@�p���c0��j�^��%�t���d��;܎[J�a�4b8*Y.f�dIu���<�n�|��<��'3�����DvR603ƽ�����X�uͧ!����"��@�a 3���ӗ�h�r� �ϑ���,�����4�����z���8huK��ˡ�m	�Y]A<��(�S��i ��,S����_A_�0vy�"�����ڝc�*���Ibȇ��$��
�bAo�0�S�O4̓�h �EL45aǨ��F4�B��^���G=��w�9�BhWKr���K��f���Eܹ��T*Gu�ԮcswG��I�U������N�=��{��[��_D�� ������G����!����-9��Ѧi���u�cD�TU4f��.'�`�b��0����K��̳t.)���;��0*���b���{Ї�}4��T��R+��c���P���ڷ�/���6"	?��B��hY�Ǫ������]DėC0<���=�x:������p�����W`��/�����~�5\�Rm�z��]|�XC0���,��Xaخ* ���7N�!T�-q�̴�FLWZ%t�$B1x=>��TZ��=�`���pFa,��˧q���a�>��W��v�gq\� ����D��)M��)��N!����He��S��,1���'���[_�#$"!�SHe���9-�G/�ϱ�yC��}��\B(�ի_�ի_A�3�j�(���Q�4I���e��VK���2���έ�/?�%<|�Ә��F���������x�͗����0�=3K[=�y����d&���̣U!#D�yc�F2��������N_��S�D
8sf��[�{�_�|�S�'�@��h���5:B*�q�#�Lg��j��Ѭ�Q'�d�XH�R�~��4�%��1 ����Z�eP<l��|�n��.TKDT�\�n�ȇ�x C�{=����7M�w�k��P)�`�.alT��im�MxdÝZ�0����_��߅;2�p�A���n���:%�`Ya��xgpP3፤�2��k�����ښJMc6
�DZ����q���R��ܹ3R�FY�ۛ��"�Nr���3�K�q]شN�)�� hh�bp�'S�����!Y�l&�G�ߣ@�4�1#�p�M� ���<Fc/j�቎�S&���S|����[����w�g���H* S�t$�.�=�{�VQ�� !�ɄK�mf[���uN���)������L�������iḝ�P������ �
x&h�Y���v9�# �$��@@6{����r��� �+��f���S	�	tL���t*����ie�ٗ��t,��M2���3�6�wv���D�m�D������R���<y�n޸�[[��q\[��X:,Y��槑$P/��NG�P�7��tX����iI�`�Pa�."�0��g�^C ��10����Ʌ$_[Y�g�Q��a���B ū��)��P,)�^�e��q��䂲�D:3�'��}����g���?�kF�ֿ��l�M�O2�h��i���!(4�w�P���+N'KR_]�qR>
x��)Ȝ=�$ҀA]A&7Fjd�Ah�y	��$�-C���N80ƶ�e�L�r��D$�3L�֐�G���h븵s�F��v��{.����#�?�9A�*����m^4�g��]���p�P/�`�����c8�H�4�a]C���)P���D������%��fbs����`
P"(K��XE�FF)����`�<m���̣��4���,.?�A,,��kM�^6��Mv2:5uI��Ec�'(a˦��i��e���&��Cq4x}~�;-�=�- ��+��s�P/�!��H��G0=��ӏ`0����h�uUl���lXa �-�%	�cMQ1�ă.�d���Eay<����N2H�sևY)`�9B��b��"|�>�֩�RR�',�Q�j{���/��krm���/��O`4�xT���:}f,�14�O�1K���쐈%g���N��F#ѝ�>�� ��e**Ls$q9.W�W��$��m��BPYmV�g��e���v��Qm�qXo�k����z��ɺ��9[y����
�?��_y_�����Gt�c7���f�#���p�?���O=�KP=�G�����W�������������Ȉ�z����������
>�c?%S��^�{��q�s�2�����%�l@Ҙ��$��Ή�kw���L&��T�������W��������U��g����k�B	l�_ǟ�?�ڻo��� ��\�8>��÷_�<>���`ia��?��?�T*�d*�����o_	��󘝺�/܏L>�W_����`>�t�Ã}����?�}����)�ʯ�&�c�n~/|�H�lD9b�������ܽ��A������
?����x��a�b�����g��; tk��Kw��W��_	�n����`<�NK��{�Nd���m���f��_mg6�=l����������Kk�{P�:�d�<^��.#�9��m��_������u��Mn�w��{��u��
��¥�1vy�Л�����H��K/~�sK������]�ݭ�0���	_4��f�Xk,qI%(�y8	��sr2/�h
�ɞ���\6j4U9C�zU��&�a�u�.\|�Ҍ���g�pm4�e�B1(lR�jf��Hj厁FO����ud���=�[�J%������=�����)$�Y�ʴ�1��i�<����> �筷ޒ�'�Wj�iL��2Н�?�5F�Q�Gi��^p��G�ia 	�ή-C�0zu`�G�V�ѫ�t����ڽ�]��@1;��~�i�cl޹.R���C���U�\�����H@���p��M�o����J# ���Y����-4�V%AC���Wh !`&Qp"�����%1�~��x��s�5���yC@y��9T��T��g��N �I�k"�2����ݝm�aO�&��d��ڸ|q�xDjky�����r��Ï����lm�C��ŵk7����F�L�;���ƶ2d2�i���Ņ�E�n�>�D��*.�Sӈ�*���6�ۺH=�K����]�b"��ML$q|绷�5��â��׫��0$�������iZ�\E�� �H�ұ���ģ	��;u��瑛����O~��������O�F���[��	%0i��ŷ��=�����$�F�ȾԱ4����ؕ��RVv�,���^�}���(2�4JGA�pvy	�s3�����A�h��c�u�1�%�ژ�*B�h#s�Yq�1�خb� ���oaj*.#�6������r�S�&�h�+�i��i`lZ�"q�5�I�u�ul	rפ��/"�-opF��Þ�1�'H27��
�yP�+�ڰ�������%#�vˀ��d�x	��BM:cC!�V�D_ȶ�Ht�:���CY�m��z�c8vöNbP�wcj��%b\��d	����L�T,H����*�ź��������χ�o	��J��4J%ܼ��;-������f!��t<.��h(
���x�lA흽��1q�:C��Ơ�C��KH���Y,�,cn>�n����`�p�+�.w�ڱ���l./0�����ǻE�gs8* �OCa}�n#È!���x��Ө�j���](� ܡz�u�P)����v$LB�6�eqe7'o��L���=3	����vFVX#q���,�ޯ�rD+�	zE�F @�i6���R�hC	�w|�����q��zG^8�E�������y�]�}�o�q�����bf�^gߺ���&�^��R����=|����)�������/|^6��~�9|��~B��ܣ>~�w[�9Y������~��n�:>����/�3������(���~��"� C�+`���3�� �6����S�"}X;w���O���'>�q���`��<�~�㟔����W���ב�E������?���D�X����X_["��z�<������,�����-Г���sO�G~�Ǡ�����j�w�턖������͛�����? ��!���~�W���(��������t��jc.�B4��g�߂�e�[���T�+�
2g>��ȋ�:2�.^�-��SEV3q�헱[�����#�a�((�[�F�z�z�b�vj��������$�Z{R�Ȥ��Ǟ���S* ������F��ɟ��Z�'�D��x�5��&��a�!T�G��6�����zS������9D��ZGu����I:eW/>����WQo�䣡��I�f*3������ǔ<El��]��G����~���|�R���xp��� ��
|�$�>�	9���y�6��������Us�XX0i�q���h�	��.�|<f�R �"��U7�/R�I�g���h2���Yi�E�0��n�L#�h�ڦ4n�I���.��KC��Cf?�H�X�J�/SX9���$�oz*�����w`�Z��N�����[��=�=5�
��Ƣb��6�ϚS��r?l��;�ץ��xDsbHؿ�U���0�d�#KG2C�5
huZ������ժ-0�����Q�RE������<$s��M`����r���'q115���M�9sF�����`y ��1V�ք�s��R��א�4��o��=��#P̉��nか�`��x�ʽ�1|w{o�sS"��ά�?����Z-L����} �/*��ww0v;H�%Q恜��nxK$�_�����菀�مb�����7��0��ܢ�������^P��1;����!���p ��pd�qk�EjjB>�18s}���C����W���(1x�xR�nml�Q4��d�sWO�����(cb:�ء�/�����'���������|�S�j���?�	��6��:qZ�p[&�� B����1���fIV�yXc�h{�f"{G� ��l[(�e����U�§�pzq�g�n4$	�X���A^K���H©�n!	#���2~ja^��G�8h��wPG"C<�9��1�W#ԅ�aW�$�[#a˼~~��&��(|.�d�9�& ������O���[�6H�S<�֘�f��Fq��wu(������z�YXx3'���=l 7u�S�h�'��K�H$OɝN׮���wޓ�I<��������)��XG0���(K��{���!�i���'�(��*;R���-}��zGj}�U�N��"��lv�S(n������H%�]n�DWn�$��0��P$ ���17Rm�r�ʼ�DJ4��St�)<4��X.2��R�]Z�O|�X�\�H/�W��o��d:�ͽ<����htʸ����?���]»�{++K8jD;E��.��/¯�$L��՛Wo�Pk"9�G[�t�����["[p�=!}��'���C��*Evp{�b���S�?Y@>�#���<��نym&e<��ihRa�ٮ��ɟ���]X@4A�VEF���K��N#�|�@��.��w��h�����7��_� �fM��� ffq|p,������6����є�}�򃲸�߽��eJ@8�O��Ï����/�|b�099���C1��f&�����}{��k��D�psIE��>,,�I"�}�J�Π/c�N�����lS�!�T�FVV/��+?*.����B�P$�`�}����nݾ�F���q��8{�<4�_���0��I��q��3��+�aww�J	�p��N�����BqO�uZ��6z�"��M��yk[z�ϭM!��`���|�����/�;��7޾�Ѕ�.އ�`��_�:�����7NE�]�j��fзg�B�4i/�V�hfaw}�1����7J�[:%>��emo��R
�����L�z��=�X�1h���^����HEx�:�a~�&��h����U����ʘa��cS��5�0T-��w��;7ބ5f4T�e�Ԁ�=�K�#�ѫT;�M�`��+L85�4�y�\r@uaz&��S���L&"���G4�F<� ������v�����w��gy.|M����ݕ���jI�dn�� Np�������$9�#!�B
����	$$�J�m���,��eW��j�����9�=Z���?��O�23������s�WA�ZCq�uR��U���H�J}B��؊R��d<m�i�fɂ�=��ٗNa9�����Z�]���K�c�|w�=���D��~�Ľ�}>��O���9,�Z��j���F��*0n�    IDATI'�����X:����8�xs^��L Ymo�鈢��r��N��X�sح��zq�̫h�J���`n�"ʅ�R��0�.��VĒ(�z�w�z�O��\HVo���u=�=�ew�$v�a����vl�y�R@����]@_O�J�^���w�+�����H��-�$���?��38v���I���׾*��}�(q�\�<|�k������pV��;�����Ӣc����lG>|�N�����&�:�t?f��19�7�߂A�@�[��zX����y�H�r��26��D,�;�m(=���5~�.�*�
��*��A,�܂��F�n_:<:3�\�W�Ab�}F�2iܸz�CPו"���G�Y���	��;v���˲65K%X�:��Zܺ����(�o�0��Y��X��\��C�W�l����餀�$�==��5��l2/
����X����f���'���_z��~�S��ܟ�ua����A��v�r�٤���h�td���mI<Xy�j�t� �6��J�R�сIG<�B.l�Rf�	;FF��,�e�SI��r�5�hUh��Ei���mb�TP���?�>��DR��MjϕDD�j�az�	���
�37%���+mӺ~��-d;��|� 4��J�l�ՈŒ"�AR���� ֹ�4�mh�%'�R�Ņx|SE�م1� �
ځAU��,./�ϫ��O��'>.8��~�K�$���o%�N}}i�0)�������7��)�;����of��PU��`��(��y�\8���o7�WPw-��$�Xe�oB,/[�4�Gd��hlCl	�6�v;����-i�ZQ�ҁ�$�
��$�E�鸒G�Z��n�R�#�g�onW�`��f$���G"��� {ǻ� q�2��D,�5K�>=�Ìϟ���e��7��cwߋ�S��'�GH���o�F��h�o=4%]6�%�HU�%Sh���`/⑸�h�(E���4�{[��)_"d#�s��йC%�"q"��[4��0�DZ�Y���UV&��E��hVnEx��dC��Ӆ�mSP�)֪I��ڱ�ֲ#��E��>h]:�ϜB+v]*��
�G
^h�~4s��S��#����E��%!�Æt:%�}$.QӋ��Ui��!-��Wf��6_�%>��0�3...J�$n>��]\�%�TD
/oD#2��HBK*���y�R�mf��l-y����V$�o�A6T�z�pTv��<�Y,پb+��'b���r(�	*.g@p.�	��	��^�5����5�D\���F"NɆTKDf��M��E�S~3�����D5��:��q}
8Q��� ��FC��K��ktR,gf��{����|�Idp�8�ɜT�z}D7"�[�Л-�&���s��0��pY��V��S�̈p<�;�?���~�R�c��RU���r`i!�]���ُph����bkסm���8%!5ڍh�k(��P4L0i@M�L��Y�#��}C��b��	���hR����0��Xߠe��5a�2"P"��l!��C�W�R�a4�z�A���>�-b�Y艞�ΑA�5��2���:��0t�	D�k(.��"%�A�2�mg�f����sB���m#����ÿ����3/��W�t��:=6bb;f0�cTG!_��������ӇD� *�S;O��͵�c�24�#B��z�`6�%�a%L�\�&��r��3g�Hatl�dBD�I�h���g��B|X]Y�R1�Î�zHb��j����H��0��;���I��n ��~��1J�S��#��@��ۄ���@߰�O�H
�J
Jpc�:�{�k|8�{�cu#
���ف�j��_�$��������;�)I�Ϟ�5�k�����Sx��!exh�5[B����q���f��-[���qP��v��#b*q��%���j5�WP����el�5�?�1����������RO���ϼ(�u#=�r�*z��Xߠ<�=C}��p֮!�������+ˀŃ��0#�]f�~�z�($s��RQ����W15�N�W��}A.\��́v����A��ĵkkعo��b�0j�|��(�J�0=>�+W�`lr��M��fLd������]���e�R����B<]�������o��_XR���|����YU'/�p�݁R�" R~��ƝqD4����"�<�o�r��pl�]�� �@����l*I
�dl����Fz#�D*�B���X=Y�*x*1UW���u�U�=���U��&5�1ste�c��GƥL��Zp�����������:e���s�A�.Z=�xj��U��0�h�0^ۖ��ׂ��uv�Lj��d�d�������c��`0[0��	K`&>��0scC̳����)W��z����;���*V�J<G>��/`%F"I=7+{�1dr!oP榍|��R�NU߉Q`�A�@jOJ����I�E� �M"���$�eL�98����M�=>N�.�ԝ�g�1�B���c�|M�w�<>�.�t
�bW>h=����^�����.@YEf{�dэ������$��%��$8q�E�/_�ˏ>��ŋ���U[<-�����/�?6�͊T.-��D�A��P�T`�ڠ�J����*+��bE����j'I��Q��c�E����fu��b�uŜm٨��OKV�l�H���j0!���R���Ѵj�~}�cP;:�v�E̟|�٢	o̥�Q���#�K���B],�r��gb��'^�����d��s����l���������H?�>ӛ|-K5���{��8�s�,r۶�I��r+�g�θ�W�f,.A��sܭ-�u-F	2d�޽[�U+�k��}�y�9�D�:k�lW�A���4�IR� ��3338tp����w��uiUq�����@�s�s�1�1�5��imـ�YA�Q��F,�-lUL��EnHi��ߏB�.J 6���#�,/��_��h7�h��C���#���L	�<�4V��Nn��Q [*![�f(]+��`�o�D0`��za��x��p��A�����Ƈ�61��g�[	�Tz�����iG�Q����d�@1-Uo�U����&�h��Y��d��*�c�����Ս�Y�7QKG��\���zf3�MMl��0��Ph��e3(R��_&-j�*�0ª� 6b|l �+�P���Z�lU�k|&�z}&��|c��V� :�ڥ��,Lf5�.��,UJ�Q�X�QI���Q���b��F ��p
k�q�-�mGL���s��J,W�-(�����
V2[���gP�<��w:��$��ݜ�S;���~[*���+;;-�RbU�l�ޞ�@z�A�d���P0�NM�T̈�}!�B&�q�� �I'�|��x!�k�~���X��F���P�����u���=���
�;FG�%f9A��D�� J�<����°��7X��D�XF�d���_��1��0�s�с册�s���V�JU[Hu�f���"��q��cՑXd�c�R�޽�1ws^�����E�v}�9�{�>��-C���jR�k)��~z�j��?B4�E[e���뫳�D�{ gϞ�Ï>��Kx�k�����S#�K���H���ͤ0v�W.�ռ�)߬)a5X�۠�)JE�L�S�H�nuh��l�od>�.���"ṋ#S.��uk	Z���j�ctp�Q������ �|lb��K�Z��A(���(6iTJuY�N�<�ݻwR5d��_��/��}�����O�����n�(��L*�w�IBĬ��.6��J�)O@����E���e��Nہ�vKDA=3�MH���T2Y�
��1J[�f4�/��`�YU�����":-�6�}��*4
5���
E��������Νۤ��(�#�� _k!_��`S�fX.[ ��⁎L�rC���6��4��V.��(����-E]��&�(�5�^ĝ	<v�،F�K<C��v{a0y���b��ch�-P9�p��u�l��H�"p�j���ʅsXYa��72�V��xQ�p���ɟ�)z��01���He4�U�c�3Aa�N*<J'0�2�@�V'-+G|�I�5БH�@�MN ��l0N��t:�Љ�{��A�Ze23�d0wz����ݡK�Vڸ;g�gŒ�����Ye�ͅ��/ X_����f����k�V�Qj�M�d�	Ga�ؐLFE�Z��W g2�t3��ѽn���������})��Ia�w{wMKU��+��#�#Bh�W��F����c�0շ$�*��h���Q������R�H�*MJ��%��Ţ#��d�Z���+Ml ���Qo���<K���x�o�*�,�gO�����b�i5rM�5re`���Z�u�xoy_���%ifK���{�����1���g�����Ʊ��(��V��I� ��nޜ��/EkY��qX)�=�q�*��q��ƥ�D�{>��0x���Ǘ�Wd�m�E6o��dl�ݻW���|=���1��|�C��w���a�I%�?ϋ��k�g��zd�s�͊��!dC=}�fR��o�"x�>��Ӄ͵+���0���C�'q��7�g�bd�D����-x���p����R�q�����o��>L��k��6�p��E<p��Z���Y��5��� Μ9�Յ�|�cx�{ރ[�g�|�zL�ǹ3?B)r;���/����	玃�΃V�*�N��N�aS�X�HK�jc�8 h��4 6/�q�Tաް��UB���y������P�Ҫ��d��>�J]!�����Uh��]��(˥�N�Zϡ�dE���
�^�A'
n����@M�^�����O��KO��Τqw����i4��E��B�C��B2[�t(���s8�2�α�I�
��͌T�9賛J�-VE����^�O�7r�1�S�M��J�>���I#��"��Y�'4���##C���E��t"�V�
	����e���dcxE����6�jH�sp�F��w��1��o�'�Cx}?|�i���f�b`�T'XJ�d�j-
قl�8��L��mPt>�L�Y��au/�g/�,���RvN�Q�/�8E����QY�d���a�ZE���Ƞls���s&[�>�'Ǐ���9�yG�2��#.L�=�N'��l:-]C
��x�n�05�œ��L�������$
��w�Q\�vw��͠��`�㡑1��5�.�V`�u��A{@6��&���2e�N֕x�.apo���?L�n�Pp �Bs�[�g�zD�V�'�=�Ê��1�N\�0��+�wm(��дp{F�Z����	|빗_���il�q^9s�(�R}]\^���Ag�zl-�����=�䟼gt���/,)<��������F[T�`�ײ�VF����(�SDY�1A�1	�[v�
����H��p{Q)D��iV�aVèS�"'ټ�\	=N�j;�-I��J-�2,��e�P*�p��Y4pu��<M#��#���䴊����1�0rǟ/V��C�4F4�(ԦJ�`�H������}��D6��~���77�ε�\����N��h�@V1q�5�jU0蔂9d�����RF�;�I�hd�ӏ��(Ph�08v����T�6��JX�Z$V7d�!������+��XAN��1\�����ꗠ3���!Mu+)�U(%)4٬e���^�f2hrb3�2ʤm�%p�U��)����e��;�Rfg���� ��L�=g`��\(H$r�q���y[t�ݔ��/
x�|O��>�Yas�'�8~��8r�N�<^TJ����nְ���ڪ�NR9�����=pym�����\�n|N3�����M������EB�R 	?A�	�r�D!�����樕�岰��"5@��V��ROKEq���L��h6[б�Z��(:=�k�&�m:���ñM�A���Э44`���`q}M����T0Z)����HR�z�)�����:�h!]գ�v!��=Ƕ�� UM�M⟸�gR�U��J�����wH�`Y��a;��dK�'�����(��$Nv���e8����qڕ�(܆#@6X<>Y��\��<⏘$��77�tu�����ޕ�Q30[q��-9>78Lj�98�y~t�)���&�|Ǜh'�8���5Rmv�y�����&��B̝z^C��v���h�PjVв���Ch�"1�?:�݋|������ah�{t6o�)��Ξ����x����|���W�h��|X��_����я~�w���~��x�W���(�x�{������<v�k6�g�x�_�m�	5,p�n�~� B��-Z���E��(:�+d�9�ʚ����4V��)h�(�5@��R�2"KQ�&�f�S��F�o�h�m�b(����_�*t(�T�i4�ʹ�f-�� ���j���@%�A>C����X�كX��у�JL�y����on�N\�ʭ�����x6j���]��j�w�իW� ��(-�B$�H�А4�m&�Y��&z{������L�H<�K�7��2�Q?�d�Z��f���9��M`��d2�Q��%�{��Z�H��km�?��贛bQG�~�Q/ګ$�HAQ�ͮܻ�b�
%��,l�~¶�]XY��,�IY�\Z؃=}0�r΄�P��f0	̥�^C����a�J����Uk�i� �.���KX��ۇb�(�L�����3)����:�PHՔ"~�l6��;�����)�h�x���Ӹ�3F�B�n���\��(�F��S��z�ҝ�z=�v��G�a5|���ǭ�6���&�@(���x�qpj��ϕ�� �\F�T����kK(���>9$�rƖV��ӧϢ��g�
�
;��B���v�f��|ˑ,���S����VT�c��iحfT�Y��1�֨���D�����z�����+_�.���>t�&��g_F��V��^Oe����r=�~Ժ=x�������?����Ф����Y�����b�C�J�"����P�*�0"����|wQ���o�	!z�_;�͵Y8�J�i>�n�Q&)��Y76"q,Ec(*U(��0�t�Lc�5�B �l�10��k6@e-�L��L�.��`�ʎ�����&��N'`�!̤��`?�2�F�B�SUiF{Z��*X�7Y�!�?/�Bl��j���-�].����ѪT`�)D{K�-�٩A��!�����a����
m��߁瞻�nL�؏K���H�°��0A���5Ԛ*�n��ы�;wI+���^���=��� 8.����/>��\�i-�s���"m���Y4�.U>��CN���Y�aY����"&����+4��`M�d��M� 2�{�z��q"q�LǇ]&qh\d����.���8���:Ejbtl�z�Qq�p9Ğ���Ō��/
ެY3��С}�6K�@�z�T��906��.$3�����ք���bea>s{�Lb��!��#R5�ۍ��of%� w����w���6"�F�
B"��|����!c��ͬ*u[�E�l01�Φ`))���P)#�J�� _WA�6���"�o��3��m�a�i�˄�p��&̖	DSj̮��wa�ժ�L���r1v;��{��5������o�����*�}KW,�;V&`������J�X��X�s���vE�s9y-�[�Xw\�%�ܪ&P��A�����/�}��޶<�qFZ�1n%�<-&�L�9v�5�rW�n+\���my��������R����0G]I��.��f>�Z�&���X��67V�k��U08�&�
�m�;vƉg^�������Co���G2���o�|���)�;�*,&�ƶ�?��(�Z]qc����>$�	|�O?�d<����>��O�7����
|����>�� f��+`h�a1�1��R�6f�b0ZG$Y�X��� ��-�c�JEB��\�Y��6�w`������lʹsϠQ�cxh��fn]A�� �j=6�6YK	i�^M�|y1��|�c�x�1{�f.^�N���\���g��'���w���"J��<��<�+b���rw�    IDAT�����U�TT�Q�Ee�>���t:]�+��������X|�R��;~�F1�@���Ng��)�'�DI���Ֆ���V��U
Q�I!�n7�%7���f:�+�k�	����6��)H�lb�Lﮮ)����{�mY;j��.b�U���M�j:
6Ym�}����$n���"�L���:��;:d�Y(Dޡ���-�?&n\cJ�����ŜX|�;j,-�šhai+a��1n��N �(y\��ad�4�Jr'Z���o�<?�VS�삖�F#fg�chhP�L���b�;>=]��DJD�9O��8���"˄���#o���?�>�sq��ī�6���g�@����Ĩw܁�����b���XX�an&�ۋB;-�xE�֡�>8��0�iB�K�9L���������{a3x��bicIƆIӃ��fn"���M����ёM�T�.]Kٕө:
��@����{��R)��'_A����=��x��e+@6Y���8�z�[C������Co����.�y�+����O�W����,�f>k���I��6 ���VE�t"`K��y�!�p �]G�ځ�>��QdWW0����sj^�*�鶊��R]J�2��9,lD%!,P����3Tt��SBA�v�	K��q����CkВUf�a�](��������d��&�=^�UJi����v6����MVA����\zn�����ixG��\h��^���A����IP��M	�@k�R���
J�5�k�f*A�7��v8�Å��+js���ā�oCN�n$0�tKl�4�&��p�b�mw�J��v;w�d�œ%�G����QԏfK%6a�lU3��M�	%���7p��	���J�$�-,'?'1��d�2a�ڹ�� ,~����_���<��"@���4�B!��E���麘�Z�ChuM�J>�C:���P������o�dP�����9�?���8/-1�;�}T|&7(�	�֩��#���Ձr6��!�n�b��?���+����c���7.]���y[�'#;X.�[�F��nWT	���e��u���3�cۆ�_�6���	��5H�2�Ѩ�����D�U�ҨJE����z� �8���V���B������&˘j��V�h
c������o�jx	:�V�9�Þ={�mʅ��	ϙ��M���?��΄��<q�hux�7Vژlv[fMy7���q�^"ԭ�&q|�j66"��`���z��ް�U2����aE�U��67��U��z���9�z���1�{��c�ek���L"����'?���g�9om���`b��PҲ��7 �bA�Mæ
��(z�����8sY�c��$��q�{������׿�-$c)�> LɎʆ{|�����q��i�JE|�� �S����7�رs��115�ň���q�U|�o>�x(���}���O@�j����;�{'&p��Kre0�oF�V���}�G�ȕ�s�����L.����� �GF�(���,��+�^Z���Ȫ��M�5�g^=�F�(��5�(w��밹���hVHG��f%3���׮������B�^~��X_	ぷ�'p�����%�t�m���04b���,Μ;�h���=�!�����~gO�@�������4Z-����]� *�xb����#�h�10���Lƻէz6�S�[�vY�j��nn���'��)��M��|��+�ğB#��>F9��}���0Q��t�R�r�����CjФ%�^/mf��&zRka�q��E�C����m�Z��6&�E8<w �DduY�G,�����ˆ�]�*���tx<��
��X�I��đ�T�
��Iaj���n-����G�Z�&��x�T�ZH���3��Gn�8���d�˵��
$�7�����5��mg����v3?c�^����:Q?2_�C���J���38u.�\Q�Ӌ\6�=;{�}j��&.\���#�qs!�+�<w��*��*�A8�V��ci�����^9���P+h�F�Á�P+�Od��6p��<T-�;4�&�Mya4hp�S������n�2��}=���wB�W���s��o���M���W������0\� ��7�����O`+$J��n�\����l�P��O����C�����<�?��|)�f�X��IĠq#����KFe:]�Bi�Za+�,i��J5��A�d�?�q��������i-8�:hZ@�P�FgE<_���d �Z١�5*4;-4d��Щ�`��|�,D�	,�W u{������b{��q�R��`3�"V������AW�0�?����Q�����w>�J9��>�WQ�Z�֘��Q�lS4���ڝ�.+zPY,(&�0��(�V�|J�¶A�V�`K<�q�D�����j�~�j{Ɛ+*0k�#���-�եeh�
1߈�%�yXX�%U+�JS�H4����Jt�n;Z�2�9U��bM���9	���2Y�R���ō���bV9a9��!)�l�v���!ck�v������GV��cҰE4�THD�t���F6�[�[�E�QH���X��j-�B6��|�<�Nf?w�_�L��ZJ������&�-t2=�h�2�y�	�2� �R�͆R=�|���'�["���^�mE�PD��©7.�g6�D��m5�&���JLV�x-�@0�0�M����mC2�����G���0%b�ȶk��iKb�7�$��.�_�X��ҭ2����_��ُ��8!��t!#���Q*X�}E�\R��a[����������U=bJ)��Djʖ,1�LY��j��n��nU���\����<���i��a��$b����y�H�``2ʘ�"{�o��:�d󼶪���*�aՂ��A�Lx�p��?�����-'%]���eB�J+���sak|�y�:
�YE"~M��E���QE'��>�ҕZ�<6�װ|�"�ڵ^�8�Ν蟸_���q��Y<p�XZI��¯~��Q,p��|�3O�~�7�ۿ�{x�/���O��g����S�v�
N_8��GK��O���x����Cx�|����y��yў�q�.�1,�����z{����¥%�k8|�i�L�V�0wc���3���Vbq�Exi@�ң��b�·q�zH6�V��e���p��*�:�/��?"�+Cc�;Sai�*���8|�q��G���N�"��^�����p���R�6k��ً���03�g�<�����ųO�3ljB9�R�U��28�4�&�ި+�0��%R�]���PEi.�R+�7_0�l:)�[��l�[�U2��М!����a�Y�'%|�Uhx|�I������uN�����-��*�B�}e�㊝5MW~�
���T�'\�>�M:!�*�������@WU�
&qw��n��F�g��r_~�i!J���T�D9ل�`G<���􎮥(�j��a���	z�^1�["��v�����r���dJ�K*�!xG!�i5��W͹��v�������{�h2R��rX�J�7_,f��<by��X�H\a��=�z�s�$�]r�ׯ�®]��(4�'��G����qr1���)��B�MOt�`W�����о=x��3�tm}C}�@4T��yl
Z�c����F"!�3�ŎK�.#�-�d���j��w�����0
J�ek��pa:e �BZ}}n��9���2�{�~���VQ�6�+F�lD������{��=sk�/]�����V�������:�+�T��YE������4�ه�������E��tA�����|Rx��������@�z
f��&����V��QhL�M0ݰڼ�Z���$�S�������G�Յ�R���ϢVàkAKW��2��"�V��Q���Z�O^�����L��ZFܾ.ˑ���
T�2�~����=�?��X�X���sH��Զ�hu��[e@��c����� �N���x镗��'� ;��FK��ѥ����%��mF�QD`�GOOb�u\8��,=�6�q�n��I�~,)_��&��R�8�5z�����I�b:�lQ4Z�j�MRk�(����X�!�YB��$����:�;H��`��G�@�Cعs��PWR�m NNJ���`�e���� *^�*+o�4Ɇf����c�q.�|>w�ܝ29b���t٧\�8	)wC' �]��lo����1MX��
T�y���QXM���ϣZM�nW���ct�NIX�Aa[/���dQ@on��0��8Y�>��d*�F��P��v`�O ��T�1�2�+���.��}nTJE�9]��ND��I&���I��?ۙL
���jY�*�Z*��x�5`6��X5�VC<�ɜ.V�Z�ly\^lF¨�H�61�c��<�=�n֐/�����b����:�y#._Y��7�	��;؇��u���9y.���t�7!݄�8�����غr��Ⱥ>����� s�?>�I=	7[-!a���h7��^�ǝW��MA\&"e�J`��k9���%��	�$񉄜/m��	��]>ϋ�G�G��M%A�8���&F�ժ���K�.I��Al�#��sz��G��
x�p�D����+�įo�T;E���?����y� v�6|�/������_Ƈ��[p8���}��&|����?�~�w~�y��ߞ�tFB+�x��G�c�6�|]R�'?�I$�1������g��'q���	/J�����ŢĿ�3X��5p{z�ҏ��ZN��TF����-�����^�}��v1�ja�}�\�*54�(����Xe1G6���l�Vo\�:�=�Z��@�P&�+-
����Ǳ����xJ*?�'�'��S��jvb�wX��N�R-)h5U{p��Ih�n��]�c5��~���)[��ޤ�Ēn'�n�*	Р���X0QׯZ���X&�j��L���j�����D2��$���:��Ȇ@��	c���̤���U-We�g�)T*e(��u�0�4Ъ)U�+z��Xc�i��lJ�X%�Y�������21dRh2wh�*+�*��6��x|����Gl�$��f�Q(�106��fJb5��Sg��i��Z*v���A/��ωj�����i;�kB��e���n�!^�婩�3q�$߰���k����é�g���De���	"��&J���B�F�Y��$�nliKw�}n(y?�����rd��y���߅J�E���|���;/�F0�;��/8|�Nq�iT���\-��{'�7&�ى^\�;�{ ��0�-BU��yܰ;u�m`a�b�;P�obqi���T��Ma��2�(^�$l?��.Q��mn@Mؖۍ��>�L�7�K��k���PFS	�
LOLcdt���	Ѣt�X�A��60��T�hB�7��[��/���O)<������(μ��j7��@�dL|��F+�-ҩ�L�Z�4 ��dq�dr@�1J�X�y�Zv]�f��Q�w����D�
j�uh�%)ۯ'˘_�#��� ����D]ѕ���U�h��ph�t{�
��jp��E�Lmܱc;��&v���w#S3��W�ŉ��#� �o�@���zx	����92�x(	�Ï�C��<N��]\�v�����J	_��Iq3<njb�OdQi��,AeT �?��xV�?��o�U���p�Ym���¨3��n"S�#U*൳3߇\I��;�`���R�׸��Fxf�g�x�.��J���x@�Dz�:��K4��t��H'3�z�j�O�Z{3 ���x,�oɐ0a��,p�ƪ"wu],�m5�Q&6��(�gUX>����������`K!W��ݖa�f�7-o��YNcˇ�l��YU���v�����B��@�A�Ao��R�|�;19yW.��`֢ ���_A4��B.�Մ�=�(�S4JD����=���?Wq�!��\�W����c���0�}T��yǤ��7�*Y���ױ2^��Iw�L��R(@�.��<L
��Lf�P%�!01H�HNQ�g�fӵ2��J$Q8�}H��h�̩�7�f� �#h+m���w��#�F*5h]	 ��$m$c���H*%������\�y>�vuk����K��n��M����l%R�����g��d$OLLH%��S�g���z ��|��Ҟ%6��݄�k��O����!��t=?�E9&�|=��e����(��E&�jW3��V$+�R��-}�s��r�ziU�JRi$C��Uo�JG� �ǂ\1#c��"_��_	+��
���o|���{;��8t��=��\�n^�S�<�ݓ{ XPi�q�]�A�5����������E�	�<s��ַ����3�~��_Ƨ?�i��>���0�y�g���G�=����n�'�w�s��:��_@�قZW��Ճ��
j��F,z3j����3*�r��Z3��71�iX-dYo"�@��E:gA�`��r�6pS��h�B�B�
���W�c=|�񋲙����ɏŅ0}׻���ͅ�O�o+dM��Ъ�
����9ӓ�q��{0{k/�F9��]�R��8����B�JV�vn��R#I���jx�f�U8p�~����#���,�`�v��Ͷ���|����,�N��5[�ť����Ң�Bc�u�)�Ut�l(�2RIȉ�?�f�R�
ZS甉�Zb��JQ�n�oh�K"F���?�P����y02�W������v^^�a=���oH�2L���gu��	A^���c���8W*JG�a�^��fw���C���h�Y-��Hr����.ѫ�+�²h���K������w	dL�釾�޲8�gŔך0!&r\��>���bo6���A|w����AhZ�)x�0w�/^����Y@��ˆr!�F�֥5�q�2݇<���j�o�f~M*�6�V�_x�,����-�7*Qln��q[a2*��)���������	8<j�~g��]LfI~��JI(��t��W��6�A��R!��*d��/a#��;�t�L���0�Fǅ���Y'����Z��d��R�7W�B�1��F&?���s
Y����t����\%7��&EI7a6jD��V3�\�dEM�Y��
V�rex=���b��e\:��mM�:������o���i���l�\�6�&B�"©"ȳRi5�Tؚn��ꈀ�Yg�İ���J�a�_�X����8mZڻ�pf�4̓����:.^x:e��>����e�u@�]�^�v�?����ߊ~�Hd�����8�gO�~����8�o��:m-.\�ž;wc9zWn�A�����0F�w��zt�,FF�2�m`��v���@�i�Ƌ+�I,�gd�^�Vq䮇��Jk�6Fj��l�R	bV3��ױ���ՙ5��G@N����,%q:-�� �Cò��j����@i�AAN>�A��P*�����s��2Yy�.���8j6���Řq��/>ο�q��A��R�	�R�s�8�L224*�������a5�fꛛ)�����g����w�8�W�JR�ƹ�c~�|� ��QX�^TU��j\��,ؤ���C8��O�N�0�ub��<p��M�!T��XZ^�I�==�I:��E%�F��A:���;KV���zȶ)�D�o��sW�]�٦ K��e�Q��l�FC�J*�J�NA\Vg�v�v�hw�N*����E*�E�X���ٱ��F[6� ./����p�Y<{�E�����@L_�R[`[$.ƒ,�j��.�j�������`�l� l��Ʊ�6q.��{ͱ���q�o:!F�B�қD��U�Gw+��n�M�R���ݖ�`r�����C*�5
�����1I�E��R���h�?|�Ɋ���|;ˀ�1�U9ݪr�C(�	��p���F�^	��B�U��zXLZL�מx�H'�\=	e}	�Zm����y<ۏ�ԙ3x���w>����B�"z�O��?2<_���D��7�����!|����#G��=�/��_������a<z߃x��g����;���G�ǎŹ��G�a��Щİo�����"<��x�̺x ���8��    IDATL�:��%�;Lj�:�٘�a�����㍗��ڦT*�8KW/��h̽8��CX����	��lv+�:�hy�Z�x�)�\|^W׮_�#��at�-^LN���V@��%�.��`in�J>�?�_�LjM���cǰ��򕳨W��ք5��e��Y$yQ�+�n�9�L�h�&a���a�}�m0�"�T,�%�a��>;'s���#�e3���U�Z�H!��l0��m}��ܢ�P)e�d���f�"�s��-[�Bz�5��4|�u3E�۬�D
������=�
2%t� &wɗxxF��\\��Z����댲���=¦��F롰�4��2.�l�2�$&�$���r���x<u�-�~n�(��k-:�⎥�R.�G��FH$�����zf�v���$_m��@���
ƆG�Jw	k\�H^�:��dj����C>W��傲Q@��E�����2�j�h�r�Y�P���؈U��K�`t���C�+������]����V#E�jL�8P�t�լD.���Y"YĹ��".��i�8��^Ηy��C��N�~͆��rʥ�����d�7����p�����v"�͈�6'�G�W4�S,J��iu���Je�1�F��Z���3��c{�|߷�c�`�����̋��tl�Z��NF��L�����R��4B)�G6�{S���}�@d��	�:�F!�2��_*��l�l�"��"ˈ�*�7�P�LB�PTKАq��6z�f�h��;Ml��č!��b~e:�N�j3��|^���sg_���Ŏ�PjL��Pt��^�e�7�@�W�jҹ�XY��ѷ}S�㯞�cq[�69!�l�#�H�Jp����Hg��Z]D��j����/����Z��r�-w��<�v+z�V��������Q�;����K�0�m
������2��+/�(�8�w���E1����E����s���GlCb�U��=y�#R���8�0&'Ą�m�'l�D��k|�A����=�?%9�Y��B��-`?-�}K�X����q�� m�vG&=[�L��d冢��q泅�`q�8������ܬ,x#��b+�;���0лMvV�J�Ђ�����-�����
�AXx�}����oE���Y�B#�ą���U���P�E�\�f*�|���,�&�ص�R:q�L#�0�|��P�Nѐ�*[r�������;m�(C�`H��J%��g)w��h5��MI0)���M=C\b%Ѧ��&��
�|�P�k���+��}��x��5\��[0�C#���5E���8�xox�yϘ��g&W��l��}��d��)>n���W�x 6�ۚ��8`eP�}�.Ə��x�=�p�N�Ȗ� }��3�8.�|�ׅ������F�ߋ���7�ǭ�2ϛcv�}���s���V�����pZǱb�D���ֆ��oK�{�D�En������\��=�q2�Й5��u�F{���{`6YX07�"gqϾQ���04q�{�����?�W�E:r�Q�J�j`����.ޒ6���-�^��C�T��-u�&��e��z��/ױ��a������4�ƕ�!��N'�!��}0*[�[m�JH�tX�4�3t'���%!"�i���NF���uK�N.	+6`Qn`bD�j���g�Ơԍa�]#�l��֐S'�;l=�%k4(�[[���Ь���5���4Cg��b�C������@�&[5I��H8l&4�d3!dSב�l���{ފv[������	7��0Z��$ջ��M:Xi��wz�`C"U��1�~��ى���������V�w�T�H�K���#�eŨ��*����@�;��Cr��EI��6�*I�Z�*|>ҙM4[q���o�"q}�{��H<!�Li/�ʸ�b蒺h�����3H7(��DKaŝ��*���Ջ2W�]�`����i����g!���DeL��c���������<��{+���s�A�I"eJ$H+Y�h,�-[㝰3��5;gw�=g�Z���]�3^{�[ɶ�`+��H�"A�� ��9wuu�x+ݺ��{�(����yx t������{��}B�Y�P"�n�!&�=�z֎��>;ѷ���Y r�c�(N�Z�.��J]�RFF����!�q��3��1�GPIR:X\s��$(F��pt+z�t�{~p�*:<�V�fawXP(1r��l9����:�V�k=�ί�	V��%"Dw؀�x��U\���͏w�?�F�.��m��Y��iA����m��!�t�զ5�K�)M�{-����BW�8p�(*���*NR� ��6Y]�YX��@
���6����}?��u�R�vh�I�r{�0�L�I�T����g~�����Z^��k�Kn������B���B.gE���?|�i����h���%@<���H�g/g���^D�Ǒ/uP�WViJg�N�}-�]��rGG[������tܷ���@K��o
ZN���d1+��v�d?92��Ņ��I�F�����Xi��;� RS(��X\�Cqg;7���:Ν?�`(���U��td��}F'��.!��G0���@$���<Q��\���X{[H �?��3sH���ŭ�%�6*�]&84}ki����À5*�ccpy�(�K���1?{;8z�>LLLI7���2�x��K�_��{�	��V��F5;�V�juIY1�:�S�o$�$a��Ý�$.vnx&�D^�9!���e*Qy �͂�'�&��L$�Eh�!D��T��n�ȸ���||���w�wHѤw��P0~�|�s�����ZdN(������m���:�Db
�N�S��7��1~p\���\���D�|	Z=�z���o������w���kE��7���UQ �<Ys�,�.��3sW���T$��fr�K�8���$���_�J/Ip�a`A�wm;�'~���
�3E��V��x�cB�n�;�{A�r���$��1��U��&54��^I��r�פ��9>
�X�q��iXx������]h���l�ި�&��髐��	W�a"�\}���s�MA�1P�*gr��'L�,
��, �>
��m��IC��olx��e$�p���'�C�O�p�K�W_�B����/4�kD��5���pT���!<_]��(a���W�!�T�,	��n0}$�B���ø��8�o[�9|�_�hZ�4u�QD"S���]ܽyv'��&�ؘ�lN�M��2T�������G���:�ǂ��P.�b�@ AgG�Q$�Q�'l��L�Y��iX݃�Q*WM����X�XE�@«��uIo�����k������G�O���a7W�ב�M"�+�Ѝ
�[��bcmv5���ه�W���ӟ���4z>ZQ̕�*���au�(;Qe�^��
fo��յ�L�����T�u�5�n���DX�WL/�y�hz�,Wd��.ds�Q����]��
����>��wo���Ӱ�|XYMct��l�QY]^���G�?��c�U-/�HT"C	�NĞ�|:�HhIE�)6P4�כКU�}�v��Bځ�I���}��i�^�ÆX���>��lz,�XУ�4��Ԁ�{�M
���?���Eă�p��vud��JE�H%�Rhߺ;���1����RD�+2%�t&���TD��@(����N��'�� @)STYlΪEy�	mz�H��C� ���q
���[�nS�o�� ���jM�y�Gf���i�m(=sb���i�`'cQ�xnV��6<>�dB{��y��@����$٫tP��4z�Z���V4�t�`�mA�����
�� &���j�J�B)��O��c!$�8�wj��m���d�׺����G��:�C��3��SC��E��&���,�<H�"Ҥ�	�F~�)��-��z�Zr~4Xt��js�յ��;�}�SC�O��[���W���m��QF�0���0�c`�x�b�U-8u�,v�|�Xr��7_�V��p�"��F�#��$�o�݆�VD$�#ѱ�:]Fh�s9%��q_DQ�v�$�
�-�w���'�{�ȕ[�[ۆ3����h0��C�Rr�[�_���Gq������ ]����Ezm��Gx�,���T<���M��Z{7t5�7��"9~��auy��@�����~��o��c.�iL$�-*�n�ᴻ�����k�_�G�T���P�X��<#���i�c'��-!�c���N~uu[�c������9+����5�]MO��ko\�7��hwDBc��U�yd췵������ַ�� �fD�oHr�x ��� <� �U�6�츀ͨ��;]���l��YQEד�Y�bZop�`Q�M��9n����]��Dr8.��"i�X��k8:=)����r{i8,�Jb���k�@Q)�*!���C�ߍŕe��[m�;ۨ��8s� o���d�	�k+a}eN:X�݇R��D,���Uj�Τ��o N���r8eL�b��G6:�U�3"���ǰ���{ÎW�x)�X�����5��8R�;D��IT<�/[�&�v�M_x�� ����W.����)dK=�=xC1�[Z��@���:��o2�M�EW_������4�>O���aE�Kk��aNԑ�>�@$����כC�7�azgǌ��h�׃nt�1J�ۖ6|L�,��?��8���[�p���;h~p����^�L�0Sz�3���'Y����m�����|����?��M?��W���hb`xH*#�L�csv�R1�jlt��k�� �8?�+׮���#�"�����^�E�`iy��Kpx�pz�(W�0Roae}Eb�67�p��q�,VT
E�Kq�Q,obp8�P4�J����z�#�9<��� �ra��0څ2��6|�q9q/��Eܚ�����sjn��˘�F��'���m�8d�nao������et��$P��P����'�
%������9���he�vi��Zkko#����'p�{�y���2��v�:=[��tC�����b���ƅ����W1r|����!3�/��'=���=�=,pTh��ހ�:�N��(��[�����b�鋿�G;���WD�Q ]���������¢:�sH&Q�Ԅ��ȵB��b�$�$��mY�,x�����bmeE��'�c{g]��l�~v��DQ�5��QD���}���R�������X�g:_DQ-�$� �ˈ`�aQ�DQ��s����Z�m 58�������p��I�f�A���4�߼-�?fXY^�����$*�#�a�Y��K��G?�G�� ���Ҥ�K�P�I����� �ə�����!�+ɳ�ގm�%cf�����T�Rp�'����}naS3)+FW�{t �ě�{3����H,���!X�s�iUa���P��ѵ��+VD���S��U8]��ކ�g�+��ci�&���ur� �NK�rN�i�&�-�C�(n=^���:c6-���Au{J��,�h���M�u��&Z��8�ؼfRIP��z`�'^����z!}�~��:=:�g�������Z^~�s_��~�f�H��R��C��(�!8�Sp�q��ylle�LI�T�nc��|��_���{��!�-n�^�v�J�7���6�Y�ɭ��el��j�j��{�ٙ�>����i��������f�a	�p��Qص��C�\���]�ԁ��<p#�ǐ-�����f%�Y×��w������MF"���`Qݘ�~]K�Z�#��\�Ad��h�T|�+ 4���C�y[�z��%��m�]�~pcI\y��x���@�є�h�����9>JwC^%�4D�ZL�F�ir���A�g��R87;vT�M�n��V6;Q��8��L8��Y0l�ə��6�O�@�s�p��1�Wě�7P3�̼��A��mM"F���d	.L��o�����9\�E�.�Ǐ��[F3챑1)��le����ݻ+Y�>������������&�v���T����\��a�>�`���+���>���1:dA�WF)G���}쾝VO!@�]�+J���4
��ZN�>�W�S�X��&�e,���OX wP���}���T�#����*l|ߙ��jB�� �"f1еm�*f��X���D.�µ�1:y'�{��n���*v)�1�� �Y�x�ns|���O��e����Ylњ��!�fP��G>y��y��$[{pP��~h����`���+h���>���_���p�6W1���,���"��}�lL<T�1�,hY�QA�N�}J7Tf*��r=���J>����16/_S�X���~h@T�|¡(
�������xe>:�|�t�4Fv�7gq��YD<��"�*gwQ)lav�&���?��^Qa	S
�dLDū$��c$�G�ń`ms����J�wJ�1�J`��AC�B(���`�������S������cn!���q�#����~G�4Hf��Q�ߧ�\���ګX�w	#��+��=�6�S<M���Z�_[1/	#є���svw7�~I� ���܀;<�O�7��M�� ���|r��k5�E�^����ď���|�G�<8s��ۛh����Is�p;�2��uIE�oK���j-/<�s8�8.�q�B	�JV&�hX�dno��6�
�����1�w���$�������y��$�|f��w��x�SQ��+���v��۸��<���lֱ�a29�+8tx
.�'OFj��f�%�uooFG�E���y�����_������/`xtD
�^��ɱi,�+��;p�%���X�F��T>�SS�Ҽ�.Ρc@�헖V$�>��:���~�S?0�F�&��VnA�p�A1\W����dB�\�>nr�5(j�@���x�\S6�L%��\��)�^s���1�>NP�OG{���५h6C�B"�Õ��bey^x��`�؀Xw)��՘U��\k�e�H#Μlfɣi"���Y�]XtM�N6�ڰڽ�N��C��{U'}�&�}&_F��Dr �^�B#���v����z�C���&)��cF�y��un��)HM�>�b�#�����!K�� ���t����Al7;�*S+S]\К�Y��}��Cw�.�����/����t�#�ZE��6UQI��?�j��^�EW�¢:���7p����y���7��
80u�Pi:8�G��B=���	���PҎ�����i�t���Ն@�N����VEƠ����8�L!��c�X���2�!�$��t<�q��Q�ugm�	2��6��E.���T�#n���*x��������^}^�NW���}m{�ol�P� 54.B�v����E8�
Z�E��#'�s37��������pw���p��8�6������@�\ElpP������uY4\LN�AOL,�OE��\$�)��VV5�4;l��=~F�ؐ��DWg�9�ڙ��IZ6������0����GC�wlH�C�בH���&Z��1�� EA_���cQ����͉���H͘�T��8v����y��IqP��L�eKmo������#S�؇����7/� �Kw�%�Bl�i��m^Jy����a����AXt����Q��zy��YB�y#b%19�D�U��NWnϢ�r�΍�����OI6o�F����e�
c)`���}DV��g���Kt����uFt�I�r��3��^����%#��&��fnq�U�������cy����)x��XX+�Ѷcva/��D�~4*U��w�:H��
O�Ѱ��'����h��(�h��G���+�(�h=�}�?�5�t�}ss��p��S�w�N�`@^K��1Fș��,�X@���X���a�P�F��nS�"*c���̃�(�*;n���:�7�ɀ��x���{͑���fA�����爐r���\z�m�H��/����������cv�*FG=��7q���bT,P�8��'�<	�M �J�*��"����n!�b�.������C��+z��7�<�&J�$ax��ܛ�?�g?�k�}��Q��'��Nay}m���� ����    IDAT��qPL��b��G�����KG��`*�|y��0j�M�����p���d��+(�:�'����~��eC��!�}��R9���!�
��,���
�²ܟ���u9�~���=ݶ�^K$�ӥ����u�]m®Tq��?��7��8π6&�L��0�"���Io�;�>%��q���� ���gps���O.\�j�8v�g��܇?"���������/��#'����ѡQ#H�ga�5��l.�\vO�+\+D�oߺ%k�k�vA����e���0s�mA�<$��V��j��j���:���&&���;&(�S�ri�&z��l��W^~]�,&*Zw`�:��"�����?���|:B����vZP0�u8��"�EW]8�hUg��bC��GOo�}O��>p
���@�N�-Q,t�0zm�>���A&}Ü��3=�Jw��2�v��iu[�B#(�"��"��g�Ql�M��6�X�t[u��~������f�F0�'�G�ہKiA��n5��a�ð�YS��!"��Pk����T�(̕��uݰ�\��IQ��\;ZQ|@�� ���;�
\@�^[��ϡ��ʨ�X^ن#ꑐ�.�J��6�,TK�^u�����ct��%E�^A�ހ���5=S�H�a���0�U}�?���q�����sM^{᳿_.��M5�pı�A�X #�gQ���M"_�"_����j".8,�n^���<�0z�m+F���@[�ڣ3���m��Ǵ���=�<�&����V�1T[� ;G�������Q��1\����|/\����7p����!�=!��:��*�j��?���'�֖7�_�x�f\R����D&k��?�GC�=��y�.����aL��1:��+7��-O�И�Ĩ�#I��o`%�A�pb�\Ajl5���P���%��'@kt�q�d��7������\	n� ��x��<j����%aՂ��9A��lN$s����bL�^�c�L��D4n���G������IcP�!�|�\��+4G��w&P�$�*|��h4~�޷	��h�������j� 		��o�&�./&F�p��(�+�嗾�X��ZF ����l�c�@-V32n;xp���b$9��Tۻ�a���P��`t}���841����A>��B��R�k��x8w� ��_�v�` ��i�����}K�:���1�T�+s�E��G���,�YT���YX3���t%3��K���Cw�������M`a�����#�J��7������/������Ԫ.��6����p�L���� "B�k�����9�g��DN��Cfǂ��S��04Qe�S7oܐf�L'�+AI1��X��$ݠ��(����}¹</�_~�����P�y�rXYM/B��Y��91��h+i\�\W�S������\�qx\��9�I}������뒸���|�\1��@*;�\:�x(��O?�@؅�Z���������Zn+[�������
9Ԋ7�~,�koA�Ѳ�*&�z���d|���|`����7���:<�.7z��C8~���&�)t�ܾ�#��:�?�f��͵U�-�#�l����C�����GM���J\�����ֆ�n��U��.�<^~���Pf���]�|��h�8y��>�|�(��̞�0t��]X]T۸r�G��̢ը�n�RU�л�ó��4�h!�b�T��4[DM\v��d-�.��5\��-��D���*��ĠuJ(׳�ى$�aU��4yO2��"��N�0r�,�vQ�Z��M˛A)�>�ݽ�^��bn���YPş��7,0��,
������U$W��a��q�r=s��Q�t�V㱾h6����Âz},ܛ�"zp0����>�3x�#��V�E*B,�5`G&[��z߸���8���E��j��H�'�U"�?}u6g ��@�[����������nܛ����<��Cp�<�|���'att8,v%H��̇?�"�_��Xc	��CP��д�1�~��5�V�lr�&R�Ǵ&��ŝ�`��>�aH�"�؟&H��8�dZ@]���Y�De����𺭸���4P��pӾ��"�T�kՠ�jȗ�p����hd`��8�Щ[��%����Ҳf�7��nN6���>��JqF��c�c	H㠒�FD���.�.���T��o×#���ԔE���C�#��Z�+n-V�^�{�<����'�X��R},��)���ZD�A$W��=v�_+�Qz���?~����_��n{�7ۭ��v�v�����%�E��`t�(�&p��ml,�ư�������O	Q�D��
O�#֫]�u���Fy��E%���%�ڮ�}�A�FEA�C��*�	5�1yx4��������s�p�^w�.���juܾ�$��-<xj
N%��!��?���4^��Q��!9���5L���p��-�"�2�n5*��t��9����1>ř�8qpV(��H���,5x�ܺ=�\�J�:��������h�jw����Rm���t��Xt����k��h�P���zv_�����
�z�:Q�������\�w����L���×�P|�f�s=Y��g���M!�y�s�0�F���wRO�L[__�ܴ�QL��rY��?�˗/�HO�e�Q��[~��+��a�S���u�T���G��5���	)X:=�JV�.�B��8�[K8<E!�"��09~��D�V�d�������-]�zG��0�Rȡ�5�%�π��K���X]��y�һ�ɀ{��A�6Ր�r��*$�ss��E3�,�9rQ�LT��܀mN�p���zω�\����)ې��f~v�ff���-cN62�vڥ#�"U���!�5���(!�!,��K�ޏ��w��#����_�� $�׷$��z�(ŗ�6M�`R"(cd�C�}����~��2��<eX���`���B��n�<~M���h5tt��9����q�
w��^ ��y`�t ��1}&�E*u*��]�[EP͕12��������������.���W���)��R����qoeF,T�ZcS�q���
UA����f#�0Š�p�y�x�:,���W�v:1}��7ga��
�A�����h����][�{�����&�;� ���ĉ���N1���6G�����	��Hy;�W�ݾ�^k�f������u�����i������Tl\F�4�bu3�^���Ex�VXl^�V<�ȇq���X\]���\�K-�o6R,�H� ���hi�\�B���c�#��\3x�ړ�R"������˔�j���ø�e�����)��jGO<��LZ�(�ӈ�̘E��Z�)��cc�B��z�b������?�P��+2
>~�4���.��U\~��Iv�;[�x�C�Ț��0�ӯ�r[����i����,��B)���� ����s'����F7o���Koab�(,��l�go!s�ԙR��"�X[)ciuW�zv��h[�;bҌ�b)�'%9�\�,�;-����3r����߇SgO��5�8ٜr����ն��v;2��է�Л����(��;����XAO5���~gƂ��T�&��в���Exw"6�1��	�Ha`ۛw��3X�{D��Ya3tX@!�J������-�tj 2E7Шg��� m!��(� .,VC�@E�F�B�X^��f�B0��{�\��jS�K���Z���F!N&Q���
X{]����
�N�DZ-T	��%e��TM3#e�D�]�5��'E��k�#�������CQ�v����K��^��/6kK�eU��S��SQ��H�L~z/�p�ݏ?����X��A��awkg��U�<����\�Ɂ��'���.^z�7�FhZa?Ǐ桧� ]i���e��]����Qzhu���<�B�@�T½�y}�M���Aq��;�n/�q���x镟�\�!�GAk`{c����cL��b Ż��v���?A���уGa(�J{�EG$vƪtDj��mC�a��P+���g�Ź''K��x��2m�P�B���l[�);�х��B�x�iY��P�6���Ï�;��!�����½y��YAٕ���t�����pq��PM�Hob7��P,�6�6yn�`���?�����H�%�Zv�,������?Oс�v����I�ȘDr~�+,��4��TSYd�g&�Л,�`ȏ��{&��J�S6�Lz��E��Ǳ##��v�i�Vved��3�ǹ��˘�H"ŵ�o���u��9}V8�<qC�V059�͆Cc#X�}W����ml��1<�B��������Y_A(���&�29�B���v55�5�)�P�6Q��D��T�j�������#ሊ+��D�\�>�Jk~��-��$ʥ���-��T�V8v�]��\X���k���PM%/7S��|?���ފf�C�_��xm�?;T�ӂ����]��|'�k(��I��(@�6�&�kh���b��}."U�n�^�l6�'�~4 7G����#C*��B�S��jxM���Kyx�wi�`"��,�/hZZ����準�2�,Ӵ�\z�Ӑ�7gS�h���E-��E�!8�4kU�:<��d��6~���01����"�{�=x�s���P��{�����o��l"5v�S�KLaa~A����!u,�͠�������:ZC���,9<1ēP�u�-l#n#1P�Y��SBتI3U�za�F������&Μ�&��V��6l�4�oi��H�X�s��ۈzh֗0}�t;.]YA���s�A`h�nG��:��(vw�2��Q���ċ�볗aU�b�^�8{�38r�All����f 6�8[:,�y?q�7<��ZA��Fzs��	��z)��\�d���O��Ҷ٥�V4�mvж���N(���$�A��>qB����{Hģ�^��<�HDbQ4[�>FB42ٴ4E4�:�t�j����T���B�j�$�<��'ˋ��η���GN��V�0s��/N�8����+����/�������|◞���	��-㧯^�~8��ם����F������Žy�;�X�}~����u3��dr�t���s���޹~���������������#(q�M���!��Iio�."a�J�2�lf{���{]��D~��ӭB5ό�5���uSmLCl�N����s�l���C)��BnYl~�m~�?�zYl�,����O�<�pl�/a 2.�'�-��X�9rb����2����@�(���KOQ�Q�b�n>��=8��zH������E_n�*�i���k�yC
9��bco�WL�m�ʉ�_z$ҥ�ޭNw��E�a��F>��x����P����/���/V+w�cR"�� 6�X^�02rV|�Ac�AjT�(d���I�� ��Df�~y�P$LYa����)�����0���p�9�����0,mT����Uxx�vۨ�s������B��ǽ{�c����;|�C��j�n��W��Md�j��JNKG����|6��f[ǣ�|hV�~�{К0\
\�A\��F�JCm��a���*hX߼�`PE�Q�3O<��O��^[w�Pֱ�:��lN����!��J�:�H��?0��t]`~v�C��}�Yk��������^�]v�6|�O����n�fu#�MI�t�Y��㒔�|��Z�L��s����0������'q3��KpT�b�ץ����"\�>B�Ѵ1�b�"��;7^����3ǖ~�:�6�\^�B�W��.���J%Qӊ����Ó��'	���؄�p��k�q�-��11~P�GA�p��|^'N;����z����Vr�uLŰ������ߺ��\�DVU��`q������y]�J���$nT+��!'�@�*h��jH@���݂b5�5�L3��$�4D���y�,����~-�5+B6c%F�P+�aSzG�qm����FKw
���o�L@S�ȔʈD�bc���` �W��Y���y�M/J�[jzQ�����DSd�J�X���������Ԑ��י�SS FJ\S|3B�!�(Օ|�x}N#Ǿ��bOAu�b����\��}*9H�z��{�oc��i������܏^�g���ѾB^��.�9d!���5�|Wڑ�{�������XT�N7��:�	�4N��D<6���}�����|Y�������S�x��"���e���ۢ�-�wҖ�#S��qF�vS����A�jT��p���G���PȀV�F-�����Tû?v~��k��na���`w�au���F��ZCC$A����b�n����Y;�֤��W�ZD�Ó�4��~X,�Y���ߐ`4*{����7���(l���Qе)�5U<���02v�K�¥��x;�F���W��D��ƃ�`e�5l�����!dV����#귢X����<1�@�놽�E�ϴ-{�2<�q,�t���b��)����b����N��"?UQ���z��Z�5����]!(}"m��`z�����Ts�2�)
���߭�/`;��b���^~Mΰ��Nb��A���M��8t�$8@��n5'�E�Z^��Hd��h�zp�mH�m�����anakkT����*=���%�Yip��'��ڔ#R��Ƚ�ƌ�wNgD�m�7~���5ER����f9Â��!z�d's�.�l�]��~�'��~Q(9ϦՔLET�)"�G�7��7�B�PWt��չ;�h6���K�9�2�
�94�iTP�d
�i��e2�6����"�Ȥ��@QkG$��I��z��a��'Ey�Og�<�h��GI��u��qtM�S������	�&���|�	>n�I(�H�A~THձq�uā@}k[�ҡ�m�%���ŉ����?�E�������U2�������{�e�ud|B�2�&�JՉpt�@�m.����9MY��Mkk(�6|�	�J�!7V�����`���9&D�>N2��Ed�ʜ��@]k��.�ir��f��������_��������?�I���p��W��g����.�P��0>�d؃���,�� �~�/�6�^��ۃ���),���㗮����nm�ը"b5��r-���2F���g?�c'�8��K?���o#T�Wj��u04<(@�^F�����4>���v����[3KC8��!�l�����0�8�_���n��2���y���������ry�c}sO��P,$#{�2é�;j�>��/
������(��9�����Aħ!��<,�u���A*�.��7�#Ds���n"|�,n�gF@�n�ح���k�'HO[�h"+���(���/!�	�0�ƹ��f�bG�������*76�W�E�tpl�jW/|au�V�[�],n��jBX����HE$G��w��qs~�;��8\�uI�!��_�!d������Q9��`�S�ׂš��/'��3�� �E$Q%���G�Dȉ"S��pTcC�M��!(u�RF<��x��u����H��.�m#Wl��![����ࡣa0�n�A"��"�4g�u矼�,���A���4�Y\'\���h��L�.��樚י��X�$�?��@��J�`[XX��_��c��^j,&��v������<���x��u4��w
E�,�LEw�#돨/߇~�#�Z�	�q�&�i<�JU�:���C�BJGC~�,���!ൡ��A����<����0�����|o��#|�/����>�r]���I<��G��z���c}u�&E`��t�|0{�\������4�������Vj�۪�ʵ�%/����g/!�cjj����N�[?x;;M�w�p{�XiD�ur�TA3�E�����?�*6V��h��ڒ��P�w�8u�)�y�}b^�k�mv�w�p�3��#��o���������2��-|�RL��    IDAT#���'q����$���8����
���ϱ�)������NV-���U���E�.���*B~;��C?_@�B�����v�gp������ā〥)h>�H�ܩ<��6�6��]��gE�L0��R6�>�x�����[3�]m
,L#k��+�/	�������P��wq��e�2Y3?|O=�.�f6�sw��	�Q�3��/>�[���=�|VD�i�GR��R�^(�M�ۉ��Y������ہ����"�(*բ�x��xX
���%���O7��x�j�^���ﾀ�#S�g��ۥ������b��x6�D��5�����蓦��b�J頋�^581�ϙ0�l��i6���O��#�b�֗�D�5k��-G�fN��E!ϥ&4���ցÓB"�Bf��:&I��+�����Nz.O��)�J��-RE��{T��zv��ņz�)�/&�P�])��̅b��a�A�w|���6嬬/zCu L���CQI�s���I��3��+\����č�S�����0���N�WJ�h��(�����s�1���L�h�8�	T�n��e16v���Yo�,K��͝6�7��ѫ�p	�M��]�v3��y�����`W��K��8D�Ë��{��ZX��A��X�n�,@'Ge��������q����c���8ֶ��ޟ���B��o`�H�sw�iV���g��3��<����"�����a}y����H��̽^���:R�(�6��uTZE�}�<t��;�x���{>�QT�~���a}��27�N���?�<�N�1�C;���|wVq��D��r{�]�E�R��w�H���S����&}���q�*��_�p����-b�l!/]'���#`r�� �6o��%S"v,�����M�)0�"��ժ�4%ۙ�9�c�0::, #H�f�d�E1!��d��NC>����� "�kJsk&s<|>zgϞ��<���]�V+�����5t{,F�����gE�Y���K��j���5Z���"��;/"n�C�o����&�!�5�]6L�&�S��Zеy�«o�ٵ"���
���^z�D�v�r�(phA���	�!$O���%����x�&<D_��͍�r�ñpO����Bd�O
�L���C���@W�pFN"Sv 9t�#�H��������A��Br�bѐ��i�F��%'��/��X1r�kch(%��R���f�΋�.�1W}�N
�EQ�wT�|<&�p�V�%AJ��ҷ�a���'R��FT��ŉ'dݐ��oX�]]���𰤭P���v�d�ʟ�c�� �@P�!�)���D���;T�s����F�)��+�T�"��j����mfR��K�0�q�^��>e�^� �Wv�����\��/��Nycp���Y��61~H���62;KpZ5�"d��䐮[�Vvm;"�(V�dᦗ֑��q�����[ӁXȀגE�]���Ӱ���\�������DE���崋	6���-�K�Z�:^��7����C��eǱT��1�g?�y���^�.���C1�<E���h�7��G�^��D̃V�c37Μz�����d3��f̚�FAY�]N�.����g����u�1���m."_/ ��w��!�4��ԋer��X٩��b��8��t5���g�_%-����4Qz�o�c"�-~�\`Y�E!U��e:�����R��` H��nǌ�[]���<.��F�L���^�p4���oêk��^�R���Ǧau:�������꘼f����Mx���(r٬�|��lODP�ݽff7�G���\��p$�sg�E-�?R��Kɴ$��l�r���>�s,��ɯ|gΜ�}�\)�ɼi/c� �d���b��YIs`��u)��w��(d��_(��"C0z��oC����"!�W9�Q2�ix�����F�"�5]��CC��Z�u��"Rl�z�������Y�3g$>�r)���^I&��!����,���������PظRx�+��p��$�˾�"��"ǽJ�}�
�b��bG|`D^g�Y�&���vG������f�`�L�t�ݫ����6|��6y�>BIT�F������'�XQ���>~.�����K������o�h2������ �`7Cr��Ę{�4
�M�x��	8� �v�^]
n"mCG�Ր1��`��"+�N�e�r�ѨV�ux@fB�j�^���tQH�n]��ã#'�\��7�"I���pY��ړ�O} +E|�O�+^���N?�_�����)\|�E�_~N��\m��!<��_����?�.�W���ñ��K����N����i@mcow{��������nWƻ��#� ��:T��rCt��H�^��{=����7P�yIB����v(����2\V��r�⧖-��^��qᐽ~�1�M�'�s�R)QZ!���(*�L�y�<�x(ssa�����Y����(4*b2����1�X�tM���ظp�x0p�ɛ�C�n���RXB���,"��rc��\s,/.	�hڷ4161!Sǎ���7kO�����e,ޛ�1C�����"^]Q�ъgw/�Ra�<u'��H:X�����4ڊ5�8t� �>&#�XӚ�Y��V���+���G����5��ˎj����h�jX�;��H@6��5�g�n�wڪ�O�6-Ud�ژ����7��N���8,;j�6�.����F�� [Ng횁_���l�"����'&ƄS�|^�=X��ry)��Q�`1�k����~cc]ֈ����<���?��c���3,��{XDR����P:=����q��y0Y ��i��{RPr�̱3�	�>���2����i2D�b򃯣�^�p_�T�T���ߊ��7>\���5���ܼ/X��y �B��31�D��u�*6�?��?��?��� �6W�V�Vvp�Ƌp(Ul�q��/A����3�mo"����A���?��N.-."���HF7�f-Ga��$&I�i�MWPӬ8z�A1RϤ�p``kK�q�*K.���[�H)8��I\�����42�~���x�O㱇�@6����Ƹ�F����{EE�~�U�n܂��CK+�O�Ү
�+���Aj�t�#ׅԉ�ޮ$�ca��u��^|�����;o@�UQkp}���C����!��I�H��l6�H8&IX��	�<H�ܨi+�z��u	@8��#`ױW��FN���ق�����&�ΘxϽ=_D��Flxn�8~��B�'l^U\,H5��D��oO|��h�w��9Ӽ{�_M�-���e߇�S���(��լ`kc�RgΞF��I؁���p4����v��Ӎ���,�����4���G?���C�,����R)ʵ#L��(H�Ue�tsf�n,���rE(�U��K�:�wRchqӿW|��(C� 6�Va�Y%����I��,�}�+Esܖ����#~,E�b5�d|,�E�x�E(?���s|6�� �,
��B�"��Ԅ)P.��~��n�@���z��&�ˁ����-4j;��3���	��J��5��^�u��V+�"�v�,�px<���B�bO�s���"���	�B�8M̉��I��r�i�*t�(����ݖÍR��I�	��S�z��M�*<�T�^_���-�M��N�*����n�!�I��������kN{��L����W�?�s�W^���]ؽ�_܎�ʑ����^��pC��p��|�DC#��VI����qRhS4X���^.��V@0`Ñi�\������H��.jv�:t�zn�7���ڨ��vazbJ��%v��rQ�p��_��������9<�ħ�[}����7s�(�,�b�af�-<��c8u�~�oˍ����"9�o��H�G��ǟ��SP*�a�ڨ�ʸy���~�<q�,�6M���<�!|��_J�HF]�8����8u�<�/{�e[v��}��s�\�r��9J݊�-!!D�d	F��k��f��x�b��X$$H�j�:�~9�{�í��s�����U��c�rÚ����������s��������B��	�����"�}#�[�;���FA+ �����4;"[�P`'YBs�C���g`�� �Cs��܎��#>3/�2cK�Q\|p�傿��ƁL��E�տ}0�o'"�eCK0a:���UU�����$6��Q)���$o ��5�)�Å�i�ZC������ceP�~��,�$4{��[ɣ#C�����n���iI�A*�.RN�7IeRɂ�C(�F���b�Q׆I�������)��%�������ψ���v��*"C�Mw��	L�B��/�e3	�8[)�� ��	?L�4Hl]��x#��h�ʬi��s��]��'Қ�e�ɔ�k�͟��`0$���'��J�Fߍxك��;2��jE|-�?��� �ʈ}	�A�I�⠧��)�`5� ���ׂU:V�4���[v2rhhTT�<��9�Z4��P��!��� @��8�6��|n�����k�?�� ��`0��ܯ��|p�dۆ���U|�l?�x?E���ϓ�~_�|>����内ߙ����(�Q�WxmR'��P,k}L�I�%079�V��?�<8�Z��������eobm�ʍ>>��?��ѣ��o�[l��alr�S�b�q��q��>1g�m�󞾁Ra�zv�85u�7�D�(V:h���>����]�zsY|�O�T�C��o�qd։��0^���S�<��Bϼx����E�R������aՎ�����7���%!яG�<��q��{?�����%�
�:V���!_���4��װy�E�6�+*ux�O���;q��u��r�*��NN_�E
�~73���E\8�]��F��m��ph:�
%L:+e�������Po��h��F{%=&ކ酻0=}��RY�T�L~򂰏�-z�YV1^�{��
g�U2��lA�@ޓ�_��r����n�$�7^I���?p,�,H�x��PJ�����@�^�v|I��u��k[��X����C3b�F�S��Q�N��{P���ꋼ�a������DG&�_��u������i"�O"�zM����ل��,&#�;�����F�%t��|���s5��}V"��K7S5�*���4Cz>g?IZ��Z�2HB�]�F�r�`|)�N[O�����=�&lf�Y�A�?9as��38��C�%+�v�[�b=���"�3��Ղ΀a���j���(��R�����dA��A ���.[�M|�&��(4����M�N������:%�}����J"+��l2�[�:t��E-M��S��Y�)FX�����xCՙ+���21�Ϳ����_���lw��0�;zJ�Y>-WkR�V�_�C�b�����j�PVc {�4���\,T�*��3blԃv++D�ǉ��p��*:Ͳ����u���1Rb��n^�@D*���E��(�յQg�#1i�x�3؎����������a�Bxx�J5J��a��b��WQ���e���8r�aX�a|���p��]��{H�EyVn�ڱ�z�n���d�JΡ��]��C#i���P�_v��qQ�k��������x
��q�/K����s���r��������6F��"^2��s�p�G����k�"S�t
��jK���������[�Ǽ�P��pp��ʅ�� ��\p9����K��1:�}1t���1O���eoy�1�V��듿�>�����fٍ�rC�8A���L&%���W151�`�����l�������"hO��{��tR�Ʈ7��훘A�_v�1��zN��$W;>��fF`7��)`.�@��s�������;[�D\^Z���auّ+h�p�)ߪ0�m-<A�	�6A�6!j�����m��R�r���G3��fI��k��������}ȶbXO�q��}�΁�+���������@U�E
Z�"w�@�@P&j��s�䚱�H������a�\��{��N���o�JrD�}����yي�Κ�'8�X�̖f0�E@�mn�_r�!`&ۯV��<O��q_���"�q��K@��.�������
$'���A�,�����u���L�����sA�+dad�����U��kw�yN�8��K�14�������N����#���H$j�Ɨ�(���Ȱ�1��t��ID"Q�Nϡ��测趲h֓p;�)q�Bh�i1��V�S=�\��i��{}�&ҩ]<��H�lc(����&o\D�g���{Y<�������t3�]"GNQ�׆�ϊQW����O|��X^93y�Th[�H��a2���~G���w�]���$���l�O����_�Fc!��{���{�q��]X�ޔ�+r�
Ţ�S��y  ��h,�B�x��}#�.�^��Ǆ^-�t!��hX<Ci��1�D�E�|��\�/����&:�l�I�G����|B2lK�<F&��lt5.����%���qv�8֝�|c�ʕ���[�r��}����&vx���Hln� ����p�Уj2Ŋ��,{������׿�B.��ɩ1s;�t5���/���OI"F�§A�V>��|�` �r�R�47Z�|}��l�������Pd�[;�i����]���W���	�-f	`��S3ӼO;������x��j_�e)#>s��W􊢪���?|�Ds2�iU��"��9+Tq�~OU��2�0�EX(�SEy,���`1�٨*�~e�8�hv�pzL�EZ+1+\��B����Uk-�=!�|n��I���څ�J�UM�SI˲X����	��nn���b� �/�vǄf�O�H��)�F��n�՟�$<��^
=��-:}C��(λ-u}|k��ҍPd
����L%[]�Ll�v�&����u=]���w�5��)�V��79wmv����a�edD#��=o���O��J��Z��F���-��4����5��n�x�\CN<�)����*A�JFx 'v���G��Sv�Y1=>�����ˬ4�J�E�ں6Fr�.V��D�i6qpbR�z\�W6��W?>1	�A�s����/<��bP�oٰ��K�I��($��v`1V�ӑ�kč�k����]�������W��3�Js�2:��6csof]�F]
�89E߆�e�ӦG3G��BK�R��_��U�bcgKk�(����&�ڧ�dfc��OLg뵎T��z�:읾��4��-��ø�����LK{�[y�M�:�Q/$VN�L9�ό�5�M�*߾�0`.����� 5���AU-TK+@��:�Ⱳ���\>�jYS�r���y�0���MO���~Z���G���c�{ˢ�� ��'ޕ�l
sS�X��D�Q��k�K��b�J���E�mڸ4���1����I��eS��%	�^. �0?:��+MU�4Y�I%`�a4��CSX_����G&_����.&���yX%���P�n�鵛&�]i�[Ǎ	�ྟ���.��
�}����J��!��DU/��ɀvϊt͇���C��6WvE�ޤ`��)�|V��$sL["(��ǀ�K�	(��4+g�~����v޲�ܲ,r8�*y��e?���ű"f�Ų\V��#mSv�;���sX��L��b��o#)z��	&5�
�.�f�V�����b��~4ǭT�o�ozމ��[*e�����αƱ��9����xoh@��)�ݸ\g�h��vr,���%n��v�r����Kȗ��{����ʅ���/#�LbxtJ"��J>{�x�����ɶW�\�JS~�I��#��-؜f�?SL�q����5V֗��k�B��#�p�mhI�x'���|�=������/~~���~�J	6+Eq'��
}�Y[���.vvoH�*�)��D��F�VáC'p���p�]�F�Lq�UL�����`�ʅ�����Qg6������/�f������k���E������u{s[گ��LO��`W    IDAT�L^�+�|ӓ�x��;�i��v	���@��ٜ�{��&S�����٣y���&�R]xG����bj�n+MT�%X�fI��E��l&�:�e~b�I �RU�猂۷*�����ʒT�3餴�ٗNđ��HE��? b7n��6���6��>�4�~�/1;��#B��o����8�I��Б�R��w�8qt�V�F.�Qx�F#U�{(���}�n�peqI�"�ہDjW*dTŒ�K_<�E)�B��z�
���G3�''��?���`4vc�\�������p:��v;�:�]]OULʠ��덝��ө��a���������`H��t\��W����N���@�s%�N�ҩ���N�3�������x�^w�S������F�p�j1�K�2е`0Ywb��o��=��F�|��mFFғ؋R��ݮz��W;վ��O�R42ұ�a����dr���+��Rf7uW�Ә��m�~�)���v:vD#S�6������q����n�
Xu�}h�9���O�k�e5���Q��=ۨ��a����[�ǿ���e��0KK%SH����YQ���A�mt՜b�o��m���	��x۠��~��*���f����B���1I�dz����ķ
���AE�w�6dq40���A�vKfCNk�Qi�P�E�V���q�%AP�j@�]Al|;�:^y�U<n'FF�4���ō�8<��-�.^1���_}�Ul��8q�.�?���-d+Y?vh��o~	Q� CA&�\�����ob1^���#8<�?���L�����E��C�Ɩ����2��F̍�<��H�\j9��I(n������Q�Ȕ
�'���Q�@%$��C��;�;(���W�	062*F������m'a�N8aFk �ˁ��q���ĚUjYJY1���[T;[;".`���z.z,wsq�ͪ9\	l�� �^k���i|-�[����L��Ί�	c#��P�@-�/l�w7f�]>���v��a��?�1H5��]�,��LJ@b�Y�����&<N
Y��U��p�Ϝ��Ԭ��R�!� �/�*���hP�����$l6��NL�1�J��S�n���%8�~؍f��]���A��_E0���-�XۖD��1�2��M�DK���r��@��"ߋ�J&�p�#y�F��7�.��,T4���HT���P�Fb�(��ʜ�>K�p{�p}��J�	XܰY�h�z�5{hL⒯�k���nOƓֆռ#�`��� 틍��c�Os���(��F��_I�&���Ūg}�]^{~_r5������1!k� �
�����qq"pۯ*�8h`/��Er�p�Jy�� ��Y%�W��afh��%i�gRi������)�Yq������D���
 �����͚W�!��mĢ!$(����¹gp��a�c w���pۙ���7�W�_ā�'$Vk/���gp��IX\:шA���t����a�Ƚ	yEQ+�P����V:���:N2G�Y��Z�eP����R�.��'���·�x�}�8{�^�jy|�5�
�6!� l��c��_�u�j�z���nL͟�W��M,^���<�~<���7ؑ�-`(4��`H��L�зQ(n��Y����Q�#���u������@:�E��F�׀�a�pl7o��X�nV=��u<������n�#w���[�����P�bh˦����B;��n�I�l;��oQ�9�:����ᘆ��F��EVT*W��.�]����i:��̹����h�ڤ�c�Ī���&9�dbk�7�^��O�V-`wo��v�cCx��122���-��?��{q���z�%�}����n��ʵ�8����C��"�����EE.��5�k��A*UCl�(��+���N�P%
��x|.4[u��갅���h��=KJ]%�ݶT�8��s�=�����0�%E�i��w��ʣ���ik�X�VJ{w��O&���N�u��
���ԑ'ҫ;'��͏��;J��b�r���k���<>6�[��������f{��`�i��-k2y���]��y9�ʜ�W�������r�i���m���Fbs��Y��d
٣�~�#�n�6{�LPh7{��֚����?�n[�ml-��������F#�s[�����љovέHY�x�mP��w~��륫��li���:L�����,*"�(�[���0�h��H0��
�7 ���<[���a J��E�p1c�ѓ�*0*�-fMd����`䌂J��Li�T�"WtQ��X�L>�ˋ�0:��?$-�) ��(��;�`ewsan� ��F�G`1�q��X�q�A��a$`E,�A1[�k׶1~�G�7������͋�0��ͱ�����"��mx�
"n�3�����B"����fij��݋>�bD����(��=*ڃ�����8.]�
��+dl.F3�(1�q`��Լ��
�J�pce]��.��*�VO@P�QC���ABq�Z{�}GNS,H�g�e?�b��ז�Q�<� 
k-�[���LϞ�S�@>�(S·�a�$D�ڨ��3���H�	\k/��D_+N�\��U��E"��K�>��9��ύ�Gf�n����pm�<�q>zgo��B�f@tc�*�F�hճ�)y�<mL�l�8Щ��k)X^O ]oCo�I��D4�Yڸ��R����D������.��Dr�M�AE��#�^-n��0X���@PHkr<I\Wh�Jr:m���7+AI7�@�-�䚘M���>604�W����F :�GZ ۫I����2u����e��j� �\x�X�#8�9c]Y\.�f�[e�9���Q���o��)� �#���s���GЖ�݊�d5�֔�7�=>��m*�9��}CiV
��KŊ�;V7b1��3Ҏ�x��[��=��9��~�5��i�캴�%b̡%�p����� �ɾLy.�G�hܡd<!��	z��O�Hy$�E(�u�GE=w^g:Ԅ;t�����l�\ś���7�r���dAl)fg��/c7��h����P�
���DbK�iuS�Ԯ`1��z��a'��jԣX�R��>t�i�iD�=��l�t��G?��=�;9�w����d�8�>�{ԇB��xL�����Ĝ���S��W�ױ���O~�S��ƑI��P/�QJ���M����P�	Y��[RmV�H����tCo1��"SJ�G��>+�z�|C���(q��������=1�}�{�fPM-ahԊT~F2�=��`RP��Q����}c�wd�3'��1<|6w��-�;��9d�{��K�������y�x�&�W�03;�p�'���1D`e��Qgz�ވZYS��d�\�cssn�+�7��q��c�frx���R��]�D�����u;0���q���+�'��W������v�y��Ei�N/@�@uQ�+؈WQ,����A|7+��F��ۂݽ8"����lS�f�:�K�M�����t��8v�ԫ��˿�w���$U]4�W��&R��N�>�x��J�X������h5�?U��*�����P��/*���g��>Z+o��\J�\�Q��b����]���{�a���R(�ww��S�z��|�cV�j�;=�행���i������ޛ��*;?[��լ"�����5����"Im���nm�7k��T���:~ۯ�����g�{��[��A����_��o����>�����L�p�q=�7�M0I�Ve�'i��}�Y-�L�H���0(5�l�*��S�.�����M��+0��P{�T����77v�UT	������\�l�bCcR������ŋo��3�?�f��M[X,�]7�n�J�F	��?����a�W*�JO��)�67^��Sx��W�s��Ǩ�,���#����D�bN{���ܣx��V�
�R���]�������D�Z��^_')'���/at�4�{�����|Cz�鄰����iw㎻��Q$M�U{��7���-R1:|Pd�6�T�U�BҦ��,�0�����Tq���5B=B�'����jk?�ۅO�� ě@Y�C�U]���v�"����ԠE����
��;$RI��F�%�#QZ3I��Iy=�Z4G����]��D�a11P>�^��������7����0w����S	
'���
y�n�+����'q���
<6*�
�{%�&J����v`|$���K��|:�d���L
��>D�D�Z���B�Z��U�b�@����]�
�R��l�n���o�ʿ��B��i�*V]Lz�����*��W�PkY��z�8��LN����r�ذVSH�SR��u �cϭ�9�R��MT2�Z�*ׂ�#Ayo�y��B EQ��u��>ᜟ�J3?g?��vC3ss�V��r��r$Y�$ e��@Zf��Y-v��,�LM	��<?��B�>ۯ������\N�ʴXds���U.�z~?�?��
�]w݅�7������
��`���+��2�Z��">h�~���h`����:�.~6=��Q�9�~4[z,߸�.����js#_�b��`����6	a}}��&s5n^�T�Q��A�X���T=�j=X<!�l!�����'�p���=�<2�%�=1��t
{=��O��'��W^<���X�;"U�r�^���ŤƊ(�Y�g���K�g�F��� �_���p��y����X8|D�ʝ��h ����o}AnrS�+94�k��D`	��ܕ$J%;)Xh��T(��|�98���ծW����8ZD£�л�9�}+�js.7NZ&��b��c��5�-e�/bt�4B�Ȕt8z�Tjd*I�`m��ȸ_Y^���H &8f0��H�2�1?rx���)����6
�����Z�N��Wnm��(�����x�Ջ8�:&gfq��w��3�Qޅ��arȋ��1���:���^#SR )&�0?5�H8�h؏R1��%���L����Y�J�hl	�����e�͌�Ǵ0EG_�[Q��,\�վ��IFFN�������O)���q�~'���M������\29�M,�����Z#�ӻ���[�ΝHd��=�����ϩ��B���'���nώ�=��x#���S�����rw>��K�^e&64�;^���)��[��&�Dg�c�ݥ_�u;ӣљ����g΃��W �lֹ�~��泉C1%�g��#z����w��� �?�?vZ����XE�ZƠg�����pA  i5{b²;'�j�!����*��2�v">�
<N3:톖k���l�j3�`d^0��=�.���v�������$�(���aL���j�;ϾLG'?q|��1q�Q�9�ݵ�����)�_��H4 y��fV�
��-�_G�����oU��k�G[�����]� �ŷ���o.ê��.lV*�
�2�V�ju���;q����������#�|z�K@�(�H|eŕY��&~�׾�x��K8r�4����v���.��+bb�ħE�����|������pQ�n"��k�N�N	3�'�eg?;v?��U�p�@�g��B�}K��X�$ק^�	� Ƞ�8߃��U&�ss����{}�ޫ(�w����-
��/l�Px���R� �ƽ�9ȍ���'��)�FGaћ��x�b[�e��<4�C������V�$���91��aP[���O@�/az��u*u�l���E+�G���j0V�x"�\��>�1jU<���H��131�J6�^���b��6�A69�&�vz�,V�,$��y p�1jH�'y�|�~{�V��?���BM��40�b�^��~������0Y�h���'�����2^�봽 hw��^t"���Jqɵ�W<g'��qL��E��rŷ�l��/VVV�������e����z��e��8<2&�B�`0 �y���Ȥ��	Kl��x��1ҒV� w�����c�>��D6�E �a�m�'�=y���mI�_����G��������I�mN�;�k��w�1r�'���)����bw?�^n��᳟�y�~�u]l����=�05b���C��፞����S�x����D2��LsE�������F�(�Z��m8�Ik�rr�Ra6Y`�y�Tu�D��D{vz��>z%dv��������5}'�~�q|��O`ei6��`T�9�㓰ڜR5e7A�1c��ҹ+�����w��>�J��с,f=u
�FOr���$r�א/mbv�Ju�:PC ��;;M�Xd[���H�p$"b#&9|�|FT�fk�jJ��?��a��QM,���{����U��^1����	�o���]���xG&�.�a�Ϣ��><����V����1�{�5�I���ǹ�p�}��᯾�5��MafvJ�I�x���2���tE`�����V,����M��.��}�S��w��/���#����'a6u`24a54Ċ�e1H,��w��ҜKX���͂��i�X���Ԫ�>��������F��趖����Lfz	j�tU�N�� ���`aW�n(P�͗��z轿�#��/��;�W�^����o�>�-�$~��~���vz둌�y�T����j�{G��M���s�{�FR�ݟ�w�cc���᎜z��>'�sa:[��L��<����M��b����[]z��v�t�js-M�f����ٖ<��m���?�C�6�����@�ۀ�5�d�	9���A�1T��X�+p7Ī��r4CG'�r~�K�TKYቐ����i��މ��������͠+�R�n���	q���h6F��k��7�P���E1�������h�ٗC�W���5lm���b��:�����uCisA��귿�Ji�8	���w`��n^��^���݂�X �|{�4�.N�����Ug��h����(��cnĎ!�A����HgSHe�h�{(T�H�{x�#�\@�^��0J��X<`�t4���������G:��v<�7����[��&�
��IMe尠PΡT)b��uڂ�
�`��q1���طF��Ŕ�߾U	�*�v��ԙl5q�Q����بL�����[ܰ�C �4��|Ph�Lڀ?$�)?�`��J;�.�ɔ��&��8}�X����y����a3�{�=-��׏���`eeU"�,&�T�:#~�,���?'��X�0��������脴}��Bg�^[�˹����h����Ʃ��ѨP.f$�H�ƈƥl�Q��vw�T����5��y���oY=�*]���<�A�[H�f�����z]�����M�|�a롪L���a}��5�k����L��K��!��F3і��x�J������󗗗��	�wM���y������k����DCXZZ��~*
+t��T/s���^[�������P�5d�w~~;�۲�C~�"�d�\�3g���~������!l��	�%�M�o�4s,�B(i �*��q���$��r,L���	Y�ⱱUM�Ӿ�Ǌ��4;�����$�*`��*-S�ݎ��Y�1�8qt��*,�֖x��~���_]���U\]>�K��l�V�Ȧ�U�dV���r�ec���6��q�Д�C�zE�-����=�g�!�j�^I�ۇF�Rڙ�~f�(~�s��l*�h8&-N�6�_`X,��:�+�����^��.�����.<p��˿�b�?�A�,f��#'`7;�����/"�]C4j���+�5R8>�̞|7�}e�B�$��1?u'�>66��c�Z���6��(���K�"::����jVdQ,.�jg^��:�V��Z�2W�*6�nU�p������R7��� :2��(��q���p]#��ܮ��bms�A�P�����x��q��A/{d�ώb��˩��ȥ�E�py\��\G&���S��v}F��������F<��
lF�b ~�c�P,�k�/"vK���ի���������yTkEd�e�앰������-R�b�Q��,�hA����lT�v���騽N��n7���Ӎ�D��t����M    IDAT�|�g����?���Bf���WW_֊�����j4zB#2�������f�z�
-]��='�Yt������l(�M%t�������k��2lwy3��+�	��}�e�����}\o��W������ҏ��:(�XDQ�vz�sf���oENIW�撗�C�������lp�Mp�4��z�
��#���� �R�-���p �.��,b�Ȗ^��D[���n�N]��cQ�rYT���Q<�L��O>���~ .�8�����-*�H��
+;Yi	fԻz4���o|�:j�o ��m����>�5�f��J*G��͆�k�64z8|؍�i��y|�K�����C�~��R	��:8�locs7��x�%���)�j��H�+��bsu#���TU8�N����Er/�f׀RӎI��mD�#�S�ew��pz�b�R�н�/Տ�
 �^��ⰟP!���N��ʄ��E���M�&d�����#G	Hx+K�۽%�"��I��5>1!�߭���!���eۏ�4e�@.���U_��p=p"A����n�߯B��ccs�V[&y��)��P���fVv�7o������~���j�AW.]����V���b��\�hh��E�{:(:�&�M!��A!��۔�>���I�x��XE��!�u����vV�� ]��5e��f��}�o�oZ��o�2�(hu[�:(P���f�	!]o���R����j5o�|�T	�V&�M���4 ^{V$Y9c����շ|���W����!<��f3�kO����Y�~y�*̪���3���@��L&���Q������ѷ�h����V�!���Ğ��F�)�.+��n�;�j�q����si4�1�s��.����7�����TIs���`NO�����Z��ѡt��F=
�>��w��"�Z�E���\�ժ����߉C��Z��6�{��p��kE�S9�<C(�먕Z0�-��Ku����R-�f7J;q�Ʋ ��0���0���8z`:]
�N��qc/SB0<���]�M��R_���Ǖ��anfJD&E�}�p��%Sp�H��؈�	���gs�0;{ ��?�Q���>$�i���{�f���d���"W�?��C�B0��S�2��-^~�����A$vN�8Hg�p����v�X��A!�Fr/�f���=���-쮼�p��\aKT�L�h�T��9�ݶ���2�/z:�}'�yL�C��E<���������Pfs��~��t�l^|*�ɾ�의��l�Ο?�����1)��T�vr�5�Ia�9�!_׀h�-޽����B(��l�ͥ+H����\���5D�>�E�X���<���1�	x�[U(=|/�{q�~�)Ć��e�g_��܉��=ޙ��׷z���{{�=�ݩ��m�F�ڱ�(F���3=�N��vZ�:����~}~nn1�Km.����W��0����񫫫晙���������f�/=��A�}�������g�������+>��h�:��bU��B.h��/�C��0�b�ZE�mG��Yg��5�fw���c{7�mz�i"I?=��^����[���0٬htT�,�m��.�6#�GbX݈c%�ES�j�N�
�=$����<lv��X�z��N��3!_-"�a+�����QW�^|٭��80��`q�j"Sae��ÅɐG��
�6f:F2�2�f�n��K8=���N�{��;��(X\����10D���I�(&}nRx�^!7ulEv�ԛ03�!�:�$^��	W`��~g�|^�����(5j��Ű�U�q�n�ƍ���墸�)c{��1���V�V����r��?��B^s��ۆ�=ǃ�i����c�0������͝u���Ӳ��}�ȇ��X&y��K+�����{p�]g��Ʊ�t��z���5=��PxD��u�/�޳N��P����8�>;��@����+�q��������ϕ�h��dF�cC��.��v1���K�o�*ʭ6��'R2�yn�{;0���j���� ���S���6+�z9����B����(�)�
�� �����bA!��/0���U�d�8~�>�\�ì:%ͥ�*�8�0بP���/Iz�#A�&��� �T�O���Cq�`H���>��
���Y�3�W�Jaew�"�o�
�����2�n��0�žb���"��g��:+|�,>��:�ᱵ�J%����C���Tds�lػ�W"�h}E�3?��V�-l���o�dkI/�2V�D��ҋO�>��8?�Z�!�e�y��M��^�)mQ�.^=���qt�9�=mL��������>���}LB���Uױ�u�.���^\  ��b�Q8,�ͣ�����"��E���o�I�X��2�(n��n���F%��ryY*|������� ��-�{O�9������L�"O3[��~�2)BMt���<A?��~��-�� ��?��Ӈ���%K�]0���UXMN�N$בڻ��G�ƀBͮC�D���ʕsH%�PjV1�p�&�z���6�p407ǀ��M8�1��D�g��}�Vo>�瘜��`hJ%��i��J��I�S�҄���ִ��z��Y�9n�F������Йlx�K�R���o���8��6�;�m�j!��H�1Y��L˥�l|^z�E�!=r�jUZǤ$ԛ5-O�n��n#���?"�������\O=�$L&GGQ�g�������}w"W؆��G D/Gf�ID_c�C���ol��\��</��ck��|b���d�ڮu��]�t��Y�+(�bT��X	����uZ��AWT�Ţ�w���w���@����	
�e��7���)�Otu-�����e��"=-	�&he$
�=�l0�\�e�p�,���pu@c 	$��Q�����)U��ȣ�l¤B~�m�AG�6�$mV�;@�kƕ�ut�}��l$&D���$�w��:�("��]G^:&X�v8%ȼ+��R��ZW��-����BU(��>��T��z�RQx?��	m�)Q7Fc{;;��#���?E�Z��m�	:5�HS*���O�W�.�TJӸ:�`j~���bc'�wkY����J���
��1��bVI6��z:�V�,lޘ�e�a��M���V�+���ǇՕLOO
��`��R Z-�}��1tў�dj�D� �I���;ݷ��R�i4096.�9�J��r��p�n�l.��@P\�\��\���I-��A��H���K9Q��U��K`lh~���}lf/<�:-�~����*)ת·��Z�_8P����FP�$1;>.JV��-F������[fz��$��0(D�A��92�r>��`mk�^�fV�0�ea��F_7���1�@�*����Ru̠�n��v�-Dv�F��6�Oj��hG��N0���N�Ѫ��26iv��ٶ�F+�x�2�Q���Q-හ�~cA���-l��M`o'% ujj;{t��KUvk{S�Ѝ�l�J!����f@�"�.�P�hqt6��!���	�$���@���
,��f4_L�I�ql�nmoH������)i��K��H��)qs��]���DBX]]-k(H���9��������lZYi�a��Y�٦惯/Jb�57� �->�bU]���y�I.5���L+���eG�iÍk�q���ҫP�F$`�U������N�$�.n�\�nb����4�G�R�F&���b�N<�����OS�n'�+��!�� ���q��Q�M�(�|ҩ�0=����2�0>=�\�������NW.��W�}ǧ|H����z�������K�ۃ7E�fÛ�Vp�Ľ���BT��_��Z���Ȟ��J�.l���;z�:����&Ɔ�hU:
G]	��C���7���w�*��x��q2�(>t��
:9�@b��$:�8u�}a�9���?;�Eo<�.����al4 3��tq0�P��򊲺�f,�k�U�$��9t�2E:f��F�v�{q����K7fW�\��K�3X��������4z�ӑQq^�G�H(���5�����A�nq*����dĥ�q��!?��~Q�<V��?#���u�}�Y\"o�T�ҍ%|��_��r�|8p`:[�ᨖ��l�ŝD���}�#�~�#�^��N���1�����w�6(|���n����I��7�Q,i�z�Iv�&��V�,��[MU�O܁��y��m@�'��J9'7M�Ӂ�bC��G>W�B��}N3�r���� ���Pm鰴GO߅٤�|ta��_�@p��z�3h���lSS�ۋ~��J^Fq��0;�09}h4����Q?+�2|��@�~|�CEJ��f�	�;�М���^��8p�m�S7�pQ�?�0�h7�ލ�K���}70�S���	�QEmP�����"�[�����h��N:�*+m)����N$47�v}������.[��ĆF��Tdan3Z�-;�n�K� +5L�9tx^�?�Xau��	�n��bl�#�Z[����V2�&*h����+zds��"\�T�����%��l!��'O��BV�X��K���)W�S2h��p��y���%����6��ChV�8rh.��W^F�M1IOv�7<.���+�B,��8�&�E�h	c���J��х9��<�y��locfnO>�]�ub#hU[v�p��A$�����ri�r]sF'�$�xg��;�O|�n^����	����M�����h�K"�i��pZ�@�--�u��d���b�K��c�b� We��l�2i�Zpc=��)�3��Q=���U\x�l���l�"�|�b�4��`/���=��F�A ���d��PT8�׮-�Q�d	�2
ߓ�A��\�����{nmm����?xp/^
�����FϪ��.�Wk�>�"������x�����d����l���M2�������,�T;��dffN�/_����8��H�q��1�ݥK�0>1*@���/�l?ONN�������;���=��z�j�ۑL�aw�ᰘ1���>��x�ɿ���řS#x�'$��`p����oGncO=��(�yok%$�q؝�NbG��ףQVaRL�5�[Ē���^A&����,�v��R�d�7�c&��iFa/! �ܫ�k���m��D��|s���H�]E�_����H�%�ܦ�	�F���3�V�p�Cx��?�bc�ڠ�~����"R7�æTP,$|��n$R��`2fE���S/�3&�!:�!�^�nl@�v�n�B�[��i��gO����~��g��Z�Zg�{g���%䗟E|�y���&�H��큛����az�6�o��n9����^��1�ÄBMA��Ct�0�݆�Y1/fś(����SF"(���U��بt�X����3���i0�Y�0������I��z��r�=Ͷ�BO� 6�{P=x?._x����=x<��e�[]����ɿ�&�:��X�[�a|f�����]=v�O�q���N��x�_���
�{ꋟS[[�ֱmQ��l�9�z:���|/U�EM8Ҭ�BN�<C�)x(�r��u{��ب�t�\��ځ\,�I8S
yU���f�^��4#[f���qcc=� n����4z�-(�8�.�=�jۀ�o����2lv�={�EM5�<�`u
@A��F)��ρh$��N�n&��������*�|'�+窮���V+��ZYHB�d0��`��;x��4��؃=ـ�d2 �$�b'u�Օs:9�p��C���p��Uki�tW�s����g?��-^��^��䤪RjX)��@l��ڜ&&=?���-LM��{h��HT���~���~�'D��b�&p�*�wH#�:����ʆ����{���?H4�Tm����l��s\8y^�Be�H��$�2��r�I%^:"�V�/��ҩ<Gk��8���َ������-C�<�r�-H��l�2ZǱ|	�"�Q/�7�Ad*�T�dk������#��+X��䟩0j����sbZI��*V�3*� �PK�&,tF��X|]	t������6/�\��τ�%�'I
Ŭr��v���N�2Mz
�����g�S��D]�'py�f���X�l�$���E�IϞD�(�׬ճ��.o�T<Iäc|z�j�D�Z���Ф��t*Go���(�]��|�A�.^��S�����)�S9�=��'Y�b�NL���z^�������B,V��p,v�rII�,��.��񑿠�wapu[�PH�ȇ�H�=a���r�n���(WZl\GW�q�_=������_�Wk��/�4�]!����R D�̲q
#(`NXfѠ�QerhM&صg�b�U�y>��k�oR'?/z���+�K%�g9\�ݣ�)y�.�����*�������A�m�vyhh@�@a���v���w�\F1�n��14@KR4_((�*�SX"5�����{�hGF6�u����V�!��P�U��4�|��'0KO�����q2��Գ�����9:��G����N*@��8v�2�T���ALVO=�cz��(dK�+�bװ����&���
��׺���� �̨������{�|j�o>�96����1�+����E��#X#�mv�V��E�&8�ү����wX��x|F,f�������7߀�7H��@o�Ȣ%[����)��$_���U�r��,���as���q�����SՅ(��D�g��p��Ff��b,/,��K�8�F�6�fK���=b�w)�E5���p���l�$�\R,{G(H�#�b�.iW��IBdfg*��}��\M$���w�ɍ'�MG� ��FnT�F����<c[�r��UN�z�7������:��)�
D�e=��)�/W���쌺G�z�Ѕ��}��$�X�>��]�t���	��5M����y�T��W(��u���^iIn����Q�j�:�O�l�������F���y�����+��@���W&��������hR mQ��R�z���Od#A��r��4��O��L�2ѣU��c75�X�'�Ҩ6�5���!]�f�Qe��\bh�U���j��9jM#�Skk�U,&;z��.��@���?�j$��>�aF�:�X���Ns���YY���dl�^x�e��-f��LU�&%ޝ�}�OL��Q�^�P�b�D��ZBbd�����8�R�j2�s?�'�J4��l��������:t���|��מŬ�ǢO���VG�`�Ӿ���bY#'ΞU!ۢ�j��T>VCS%���c�^:���������x���w8~�0��N:��\�`��T�����+2+�<I�֥\)(fW6`a�D?&`P��ץ�׮ ��㠩4D�S�&)�Q��H�\��p��ho�p�T ��0�L6�\C�ͩ�����@r�ԚF�Zemm�@�GQ���ިb�`�3����)��,�N�g�&��*s����7���=7r������c�}����r�[��9ǥ˿BW[��\!l3�1;�
����f4OE�qi���;w��&�O��L/�c�x�k W�as��[L�����!ń7K5�W�Y�a6����M�SRt���Q,��¬�F0����ռ�#�כ����S��1��v��
l'��Dӎ�v�`�A��[���9}��|�_�8�O���5�[�}�,���ty��4�k�Fd�_�US"�J�w���P̙�~_@BdD+zOY��=
�ٌ��Tp�ץ�����Y�+(�A2���`�rJ���0�+p*zMh��I���>q0��T!�Yoi�e��Dcj�+�W�XH���˕��w�����.�+q̋�_@� �͛7+9�2��� %�V�NI��ŉ-�[��y}��L�R1���d#S`�M��NW�b���Y*��t�� Z$Qа���`l��ܩ_P��ʚ�cǮ16v��Mc8�6N�=�_�����*%i{�S��yE*11�##w9T�Mf�������Μx�������5"5)���҉������j�(�C}=�IwZ�Q��wHq@���I��<�b�lC�gp'u[n�f�Y3������'�QOx    IDAT�,cy����i����M%��%��c��Cc���b��)�^$�>I����oYZ"M�g�>��8~��\1NN���֍�7�'4Lw{��iN<��Yڻ�� ����=��r�)P�I��$��ι�J{�78��F+�&��Z�L���a%9q9�J(�����{�p��)������7]���Da�%�M2�d}�!v=Q���$��6�P~�g?�ܙ�J�$�y���=Vb��V�9��1�&�F��g<��[\'/n�p��k�6@9Q�r9P��m�Si(ͯn�u�=��y����������KK�,�����������Ժb
�5��A�N:�S�"� d�JUs��`S7�d*�P����";��a��Y�[������vI ��F�QV��ĩ)bq飵HeW�ICcd#�$R(-�Kl�d�k���*V�m{fva�^�	���B���<.���w`��n%�ɱ{�n�����E�˚�^�Q�4��P69�mDW1�m5.�U�8�45E֗�r��_`����-5p�صw���<��5�f-w��*��Xa�՟bl\�eMR̥0Y�,D�ݏ��n�U'SK�(��^'�uum��'ߧ���mC���[F����Z,��3gy�;�R!�f\XL6�z%N�z�~on9e�K�b��ʵ͞294k���|+�C�m���Y%�����h�3V�#W̩��j2��Y4s�LJ$�CǠN�F��yje律F���7���$�P,�|����y0(���I���ng������٦D�F]���9VW��&�&��΁nQZ�d<�^��,۩�kd��$Ǟ�:��z����sbi��b�|���l`����PX�����������c_� �Z�UO&���ԫ���l���},^^���g���~�-�ID��Q��B	O8����d�[�Hh#�T-4v�����9��v�Z]���a�&�k���I�������x9u��҆���M��K�9z��s�Xm.,F�b'����s���K�����*�u��Z�A�1�GR��4�}$���bP %���#�Ƣ��{� =�y��*�7;;�7Y3�m���j%��:�ډF7 �C���r8Si�ꭖ�ӥ~�4�^[��C+�W��8#�ހ�ao�-��EE��Z�fU��T@
�0(,��f��!V�<�����X�=N��h��:I$��MՍ.�*��{�:�5f��kZg��/����{	n���d�|n�K���߷�tFCS�Ↄ7auZ������s��m���z���O��9z����ʗ_y�\���w݁զ�G?������o)����E^��SXty�����:�ۯ���.���<�����|��f�k�BYb���Ke�ʗ6�eV��&�����4��Iz�������yΝ:�o~�c��l����HH*xV�*a�6�-��LR(.(�[�������I!���s?%[`�ͻ�Y��밣�j06,,Oͳ}h�C�|r�h1˹�ں����glL_�¯�E!1N[�4*���$�8��T�Ա9dRz�q���z�������9}�F����[��S��hw�JeX^ZQQVG���α�r��7��#�v��RkV��jW�Qa�%�*�J��7�=����.�xee�����͛��;��$>��Çn��/��*����Z���{�g��P�C$2��.��E����Fg�X5R�x^8r���l�s���Bo���+�A���?�m!3�~��N�VP��Z��n����Hn�rSu�}��m*<3ݓ��/뫋J��uZqؚt���<8̥3�p��|nt�
���:�^�ȫ���:v��5�hf"�*����J��	�u�c���=|�țX�[���{|�S���0�S����?g��[8x�>.^�`�@�g�/����=�FL�d�4�N?����`���e<V��N�V+��㗏��SO�Z8r��T�&n�鰺&���޿~�����d���![e��K���hkr=����f {�C;o!�����fA'�Ŵ���|�t"�������J�����ߞ�O���2��i1?�D����R�h458�bO�f�Eu���6�fZ.+FE��^
;#/�/,�QoT��`��p�(�L�PPm�Z @�z��<�dS�!z>��,��`�M�>�J���Y���f��҅|���^�[wm���!wH�R���Kج:L����VV��v��;���*��Օ|� F��6G)u���	j��\�v��t
\Nk�t�}�7�\YU�Ӊ�:��F]��ML���Mtu����1��� A��s/����e�VN�|��Wρ};��l,o`����lԵ5e�)2*w.'��R��m(�r�X��	�;��dn�*n���{YY_a)^"�0�bR�a�p?庅S�gј�ld��ِ��),��e��==��}FM���8�m*�D�]r��h"�G����~R��2�,./����bU��e�*�~��3j|,�PF����r�p&_�>(�C� <a��Dt=|Z�U�m��h�U����-_N�S�����h�EC�U��Z�W^��n@���
�M��j�!S9����6�8�xB1~�n �M\^������$�_����"3��ۅ�jk�~Wk�u�Q��YĬ]fS��&K� ����<�ͯ��Ķ�[8v�
���;��֨p��Y���ws߽r�;8x�m|���U��7?� �Ї�<���{�����}��ė��e6�m��˜8�<.���F.���Z`y}�R���?��|����f��۸z�'�LQk��B�)�:�h�b֥���z�8�|���z�[�U���g����ص�=��f¤�`5h�5*�E<Ni�9�ϫe~j��M��a����E��Hj\����If�l���7��;����D3N_�@�n�#�.���+��ʩg0�dz�S�]F�F�#�A:'�yZՒ�j�ͅK
E�n���klĢԤ2P����:�)�Ew�����FyL��6I+T���;Z&�Y9�-N�jj�e8Y[^�e-}���ϫȤD6M:�a���nV�V9\�<~B��vf�|�f�����l7����v��ï�(��"v���J�nF�?}�η?޻y��zt��x]W�u�ɯ}9�����N:U��rS��o�V�R�a�Y�hģ�9���被c�b��yq׭�����W_��,�;Д�ڷ�z!�X&CY�|פSE���̠�'"з4
�d
0�e-����=v�n��s���o���<����{)W�\�4���
:��}7݅��Q)��8�_}��<N�Z�����Mΰ{�Vg�V���"����{�PW=,�^�����#�v�.�|�mҭ��s��ʕ��q���; Yd��/іO�4��굤2P�t���$�Z;fw;6����e2�yY��b}cY�-�����=���*�K������s���_�\i
ۃ���Vh.C:�`x�&��,�߲�2V���V������5������	8h�
bʉ+��D��&/�{�>mmU���6o!�L)SPN��Z�u%]�f�-���e5!�Sуɺiş4Ժ�Ѫ,�����B�<.FFp�	w328DdE2��8\0;���+J�m�:0m��A�m]�v�r�K�Nt}�ဆ��4YX����*]��,,.�w��� �xTU��9�E֙^\a�H7��(��RYM7��CK��F_���i�=7M��a�Pkd�U�p�+�%̶ 6W�ɹx���9t��lS�!�Z�@0�\4���zIt�1�f6���L$���L�B��ɋkd�F� s��&D�iQ�G5�t6�V�� N�\���'�j2��# _����&�b��A#�b�d4&��_�w��V��ѫķȚ��SL���dm�>U���l�v�F��kϠ�تVۂ�r��D?d����z���C{j��N+0(�M�ݢ�ײ ��zWa�-��-�!��XqG�(���X�hZ�����dl��W��V q�.zm���2��
�>�'N��c▛FY�>���ɽ��	���|鳟��H�6��v����}�鞻)U?}�?��Ghh���|�3������x|���������/}�HE�|����K�����}��si���b�ΐ�Xd�@��ʆdwjx職�mX��4�=u�Յ>��r<z��>�}���,�F�\)Fdm�N����{���׾�u�����>ĳψѫ���5
ٔj�r��XM�fv�L��e�O�̸B>���x�Z��d�{od��K���G�<�k.�=���gt���a�"��4���U�z�jɪ[&�����h�T�P(XY/c�u�9wiR�.��ܔï��W�Z�����b���J��5���SdM��|�F ����Z���a��%ҩ��.��8��4�:����u�aڻ:�$6��3�!��=��u���ik����`^�|��<�(��}V��+�29q�Hj�p��`G�d���w��n��.D������~߲2����%�?h�VU��T���AEψAĤ%_�b�z����Ø�m�!,V�/���2�a�P�E78��o�:,�UF����"#*#�&�j��U�b)�*��&ow�U��l$�J<��l���+�x��-objb����
�<E�5��xU���wT_�դ���W��?�5��ShM6%�p�f����ҸIl�z,�;��>���� r��W/�o��B�&�^ӤS)��4\��mr�5n9�07��ĸ�ʏ1q	�=���ͦ���c��{�&�h1�L'X_������S��u�\����K'��o�H,Wk$�d]C�f��
���J�5��Ӡ6C����UcO��P1-�V���R�-����H ��|�b����R���]��
���ǩ"o$�NL.JGXo* �&﹌{�*��{Zyu���
����Z��F��
�����R)q;����=�6������`b��:PHL��,L��Y[�7���E�����y���ؤI$�ɢ,�j��cx���n�2�L�X6�R<B�V�������`sr���ӹ�؍dK8&VΞ!��&�����t����-n0��N0Hfs0D|y�Źq,����Z����X56R�������1b���w�I%���-Ƙ]�`vt��R����bq]@�8�'�ђT�u� �[���r�	+��5� i�/\�)��T�o�&�Y�Ø�~���& .O�ϣ���%�O@UtcC5jdD4�J)p(�+�^�n5���:��ϙ�a���X6H�Ps���&�F-zX��3�M��"�[�d�գ�*�v]]��Ri%E��I�Y)����"��X�կ,�+�A��b#M&���!/�H��&��n�����<ck�a�B���pR%M��F��R���{�~����)f���Ma����駧����s�y�o}�_9}�oy�����x����/���}����p��
��g����U��|��G���8s�4G_}��Ɩ�>��.`�D)Wc�
��G�o����I�8��fU"����,n��z]Cti��]]*,s{�g��p��;������g>�zb�[o����(m�0��s��U|^;��+��q��	z��yK*�v��d���ܲ���>�_�L<������oV-=~���@��F">���iŤ:�������Q"�'�������c��N���NSrE���I�����+����:���
џY�-�	�%0��ʢb�� !����J��j%9@�斊jtl2�Z���-��sؽw�|���*��L��g���aw���ʊ4��d
i��}�s56:���.Ν�Z+���R��T\Z������#����=������h����
�.P�\:fy�����bn�m��3�[}�����0]��LA���M*�à�`m=G[����.N�z��g�������&n���x����Dl�2aO��.>��j���e��d�P�g-��L���r�d�A2�!_��o�m7Y�r��Q��x+�.%�jLL^<���fn��ff	z�����w���>������U�:�W�S�6�x>�N���y�;ߍNt~�<��9~������X����+lݴ���sxC+��}��{9|�c��䱟R�'�+�i��9�0>�`�da9��lz��B�� ���
V�9��,/��OdZ�1�y��.fW��%x���n
�Y\�Sfq[�MU���*��J􍴓��N��׫� Hc� GaE{f0�In�T����
#'��M�����`O�j������S�����z�>�b������/���r��f�l����\
@��� y͢�X_������oeei��~�}b�y̦*m���.L���l�hgjz�Z=��k��6b2���s��2IV����ȡ�=Բ9��U�6=�/���u*&J���P����,&<�Q��C45^4Z	$�0��r1��.(�IG�X�LLNcu{�&'���ѢF��^�a_�xt�ǁ�l�/<H��~��#m�����&���(R\�]VuV��c�LI�q'C�(4�44n�V�\�p��H$��E�����[�Y��P����a׮]�5��{ѓ�{�l��e��� �b�O���L��Æ�K�C�q��� ő{=�H�ɕ�X����&c+]^��W�U����֡Bd�w"}�TK���;��!%�eH՞Ā,,ε�qt��(����
U���ݡ�%�s�!QC��bsZ�E�;��A>W��#����C��u�VV*�T�T�y|��S�l]A��t�&�Z��Sǘ�9��X������/Y\L���ǹ�gx�����|�S��qӭ��Ȓ_��y����/�����/���}�������?ţoy�O}���,���O~��z��~�OU��g?�i����L�y��g�Tˌ_���P�%��z��[8w9BW�~ƶVQ5��^���Dí����hZqZ����/��'��y�w��1�ڷ�A�0w��I�#��v
�,&� h�\���R)����v�,�=�� 'N�P����69�K%�,.-�7����FGƔ��գP�`�l���ȾCp��7�X?���Q��560it4
���!Bc�|��.�R_��^:CW�(�XA��D*O�P���e)ˁ�i"S�`���h�,,oPo�i�uԛ�`#���D�(L���$�V�H���|�ۭ�d�P���R�I6i��v�|����t<��f�R�qr�z3��k�FQ���xD�_�yI���\Oqq��6	&�tn�᡻�����e����W���
�nPx�����Bv�=&}�|!���5JU=պ�R�N�X�M��0j���p���cʠ"��R�������n���w���o"���20��m1P���%cL�~��e�%��rY4��3w�D��B$��|�g��|�g+��s��N0��m����Rrm�ή}���?@.�diq�O���1� :,�2�H��^�QSc��F���}��}~��o�N	��������WiPd��*rR5���)f1['1���p�c�y�|�K'��h���̑ɬ��reW�hMm��ML&+�T�ZՄ����039=O!Se��V���t�<�vm��������5�<��n��RR�#�&��t<����}�^�&��l�2�Sȥ�:I�KFg
��W�1"���8g�iTY^YTz���0�]j3�.�l>���|=#nYq(
c��ݫ�c<�V�%���dJH���z��4��+�jfj���.5���i9�h�d��bsx=&�V#���i�֤��H(�&���,������9z;�U��8% �����{Y�8�A�%[����c�m&�� �rಹ�22�Ą�)���nڇ�1���T\��-\�0��ng�P?эU�I�=}���,N%��<�@'�^~��'�ڪ��F����6ă��W�~j�,����1b�U�M	o��0'��5n��-t��>^;~��~�3\vټ�Qjk*��n���A�q����hV������X4�X6aLͦ���/�Jք0ɪ3�&̲����ZC:݋&�$�!�Z���)M`�����&��E2���`ll�ݡ�
e�U�T�A}�*3[��Hբg��}��k�>��^�(@U�W��R�  �@a��0��V��\�ψVR/�_    IDAT�^L,�p*�Z���k�����R�L2�S����m�t`��r~���y�G_�el�����|������/2=1��;�cm-���y�G�N�W��]�}w�}������Mf8�#�<�'>��\���O<A-S�����������'��q��1V�fq������N"����=󃧏2�P���uky���р'�e|rQ�����.3�8��e.��1G��2����Rp���?����_� �ݬb��z��Jj}�Y��ג�Ƙ�t���_q�S����yW&2�A�W�L-̨����r��.�_5/�,N��x�G_��������C�Б{���e}�8:m�z#��ZU������$��bT��j���#��X^�S�hp�<$RY�	�a7�"�h"��d!W�c�x����N�6/�DNť�Ki��w�u��vY�@��Ț�uͪ�f�=N�oi�Jl�غi���4$(�S��mccY�]V�A�Z�UC��U�peu�`{@e��jf��Q���J���@{_'���~�o���5���c4���q���u|����:}��P�N�S@�b
�∕�cM��|�I:g ܽ�F�N��v����A1���WT�B�`6��Z8�;v��oǏ}�rn�z���h�
,��au9hH�`F����}me��6��'
Z&���.�x�[����[@k��8z��[�y嚞�'�3�7��n�Yר�� ��7�F<A]�Sy��B���E�J�+u2�"�>�>��Q�KSA�l6ʷ��u�.�Ã��wPiK~����h�Y����7�d�L}�j�*>_�tv�X:ΌĜ�:�ƅ�k#�뢽c �-H�� �O`s��:�<��g��/�.h)�sK�`�\�Q���*�
��+�&d��a���7�z]m油ɦ,̜ă ��:���Կ]�m�3��g�	�˥jפD�������&.`@6�Z��K�\R�#n[9I��P[���Zd|'�'cAѥ��6�:D�-�%����ؾ�T|��?WǏ�ld��J�����Y���m�ý,,�(�f��auu�Db����R&Ng��f]r��6:Į-����㶻���a9�䰒.���va�)$Kd�i�Z%�70��@���3�J�����ի���]<��K�7;]N`�;)�,,l�d˖�x\���,������7K�R����҄�#~�ø;�y���7���6s�Wh��Rk�mj�[��:����-~��,.�0j�|�s_��ͦ�V*�$[,��|SF�5LF3�G�A�٨4xKK�
<I���C��h�`l��Rɦ�I�o2J��I4|r���$�L*����jS�Kt�r=lʿK�0�R�' M"j�9.&�	'R�����@t��K�^���a�|
@��p'�W�7yM�f�ϭ���
�u)�U^���T��ë�S L@���*�SoP�-�! ����u�*�6�|D�Qu�y�;~��ێ�a��ŗ��.�{[��"kYn{�O�h=<��o��O�����N��#�bt��jM�>��O�y�������"K��={�/|�<��/y���y�F�����h�8r������c|�*/��,�j��D�%��@j���C�����<��s|����������ի�}�;v�_O�/�hV
�����)��Cw��ޭ��'�It=��ߧ�/@2�A1[�%9�*�چ�j���˯e�ꋴ;��26��Μ]$��'�)1�k�������p�<��0���R(��4�x�_��'0Jvf�~��ַQ�;���	t��R���ٝJ�#?���	N6<	�/VkT�.�dc=���u���b����%�Zt��S�X-.J�:��R]��u��lA�`e<>?�jSe��VUrRE#��%�{]���+��խ*G�>��	�AO9]���s�xZ4�.R�:�V�Uh{[-��ĢZ:��H\����o����hd����>[�?��x��p��w���N�Mr��e��2R(�ɦ�T�.��h�+L� �+Q����Tz~{W���>��N��9����C"3�O��+l�o'`���=�k-�E���S�W�[����p��Ct�,�j�َ��%��pe�Į�oax�=D�1~�VM�o�_����.����c;�/ �ʕi���!�������|N�6���>�rA�9�?w���DWO��W�2�0���2�;����A�'��˟<Eg@Oo{�j�����C�݅�:Wν�A��^�"���Փ��X=�3�6��̝lc��[��]�$z+]�t.�4{��*�B���0�Ο�\50��c�چ�ii�`7��P��XU��B��I<�R��n[a[�{�ފ�P�~�F��1��*�9
�#�C�lQem)��V�\-)  �_��N�Ce�	c#`D4��A(�X���bU��.,#k�˦/!�����%>D^g>�Q�@ �T�I�E8�'�wE��&���fQ�?H�ž7��5���c[G�⩧��J9�M4gS8M5��47��mת*Cq�&$Bey���n�.���i{:�C~��5<.m�f�W����F�lԱڻp�{XX�s�#���O�7�I��V����lٱ�;ҬXx��Q����n��i�2}����)��<��Oлy/����}�]z�V�K�����<\����0�z�{�HE*<��ϩ���)kQq�z�iH\����&�K<�Ҕ�F�2���:ek5Ri	����y��U���?��G�\�ڒj<�aɎ|=�F��[!�A377��d,���Ȏ;�ZײtG+p&�Bq=G"�a���={��<Aa�e��aF���&����/�'�<����j��-kJ��E�(�U^�u����e-�.��r������S�
���-�UN�d>����r3��r�&��2K�Sel���h��C�!��r��I���/1�y��T�][�v(�/�)_��o������Q��0_��7�g���~/����8y�5��~B� ��O_Q1@�����'�Ϟ�>��
!��Ht��@�^���mo{?��y꧿���\��y��� �|�B���a����1x�%7T]��>I%�+��{�˷����?P�������O�	F{w'�b��Zm�Ɉ�V'�q�y���0��},�Wx�'/��9D��&�f'�R��M�=�ųg�~�ή�uΜ�9�/�oV�r+o}�12'�.�A'�cM�f���h���S�i�ʠ���h���^^>y�B]M�&�6�6�]_w���U �h��Wȗ)*x]�$�Ʈj�<�RU9�ۮ��s`7�A��٠���d��k�ؕ�Ft�"CpY��<��	�Y"�K�����Z�㲛p�-J[-U�c;�������Sh-u��^\�]O{�u���o��7�����)��������� �6h�#���%�5�+���wd�	
e9uV0�$��k���4�Ki��W���u����'����p�.����%n������T\�/��������2�c��MꃚTk�1�I��L�j��`�8���5~��ߓɬ�r0�F2S=ʉ�6Vb�l'�;��7Ҹ}"��)�R�X�f��ȃM]mܰ+�kS\����豗��n��_:)K$�װi˄|uj�#�尿����s�����fU�I�68zf����l�|'^�H{g��t!��5Mm��}�[l����(g�BIN�=_���t��B��K!��&=��&z��۫�3�� [#3�b�D����U�Iʆ/�O���
xT!�6�|���V,��[ ��F��_���M��}�*���r�T��ժ�2��2Y��e�(���=��z����(�t��ٟ�c[�P)�1IX�E6��,,���_��7?�({����Ԝ�4�r��dL��`�K�s'�^㵗��M^<�:�&�&�8;C[߀�"��CUc�8q��,,�*�d��NE���*f���u��7��	�1�}��(/?��reڤ��.��S�+<��w��7q�k�=w�c�^��;���x��E��.v��^�n�<��W��QĤ���,�ժ���b)���d�ᱛ�����gp�\D#��&��aWWБ�B �\��z\]�ޞUM'�(�@w��e&�b�W�&T�@*�P�����z��|��E$�I_��ZF���r�Ș*&�Q�����E�(�|�',����x�f�fU�J[8Ȯ];x��'�z��T�dt-kV��z�Z�2�����7�H�P��W�*+�I~y�JU�{��~�x<ي���q�<�y-r�J%�*V����x|���9���/�H_gc�D|�w��COXG��LM�b��w�n�_<�4�<�3&�M��3��]��@�&���'������At��⋞-�L�wY��Ll,���VZ7��l�:�B�C�®�3u�
�6'�z�ZS����ѡm���y���yӛ߅�k����`h���V��r-K9����W.�ji���+��'�o���t���/>��Z�n�	_��5�p�������E�[@�����q�2�{c�5�}--��7�pپ�6�z;����F�Ѥaen�A�f��z!���9V�~�YS`dx��짴0�:	:�jR)O��z�0��׽F���8���%��u/��o(ǲ$X�f%M�.sH$���T)W[�^W���}#�6/�RjjY�ĉf��\�ڂ�;Ts��5�&e4�aX�׫����*��++3a�P���P�h�^�P��"t�=��j�Uh�Y���,%�0:�RU�zn{j϶����S�z��?�z������&�}����[.�x#^�U��W�	+��~�#;v�gu9I:�&�R��1!7�e4:#�l���Ae��0~�l3Ϧ=��y�'h(0�42��asr��8S�4]����|,�M��׫@OiCQ�Ec �i�1r;��ī�h�F~���1s�=�=j,���<O#�Ūw(@�;r���qN�W�&��z���_ҹ<��l'I)wݶ�z;=�L�c~�>��G�5LN#f�I�la������a��t����Z���+h�	��*��Y:��(V��p�"� �� k7���dl�,���۷N���^Pm���UNLa�͢T���3�+�AZK\� &��pSh�Z�:;��bJG�*�D���*0(q��/�#��[5s�a
�$���	*����j+�()����\h��mf�r�@ЧF��J�\6K�\k��e�JVjuu�#�
�.W�$:3��=n�b�$@\@HwO'����U�k6�"��L<�J���T�)����;���H%��0��x�v���#4�Z���\����ˋ��'�5�,��)�T�F�v[+6%��.�R]���i M�KJ�I��@�I�� ���r���(�h��'�3?u��H��C�3Qӛ;p��{n -����21�-c��*�%��J����m`p��z����i�[Y��$�(G�8�0g��X�C�\�fh��4ʢ����e�t�E���9�{����ʢ�h�XV�C���l6+3I[�K�6y�e,l� 6�>y�dM�:��U�g+��U�(Aԝ]*�M����	8������12N����'�N����aLF#�N�T`MZ!b1�A���^\�Qս-��R���I��K�Tu�²:������~/q�S(�뢟���ŅU%s�X#I�lFe|��4�ӢG2&��
�5i�����c�i�u�Z�#���7��˵K��g?�Z}dd!�tl���<��ٹs��r��O��َ�nR5��D�̈́��Š�l�G�t���u`qj���~��&�45j���\����{�K�����O1=9�-�E�=Ț��H�K� �5��a��m�(��V%�q����yۃ7R/7y��9�U3G�<�?&��)�����f�I$1Dj�s���� ��b1��\Dce�}�{��P�&&� ��A��%��R-��5cL_z�Z~�vmf�͋)����PN\�^�!2穡�7�+]b���������z4C�X�n5�����^���p ��L1�W�
ʀgw�/�Z9�J8�Vb�$O���`����$se:{Ued"��v06�M%�DG�E�@�0��fck*"�L�Z59
��Z���$&C'6��^�۪�QHb6���Ag�c���\����S�|���m���7��o��{^S��`�z�+�,d����|�?񈀂n|�A��U���Hw��1D)�����ON��� ���Hjq����z���E�oo����4=��}>7�Bo���������J!N��B)�����8��5dJ��N���t�x��g_�駾H�_�._Q��s��:��j��d�f�6�V��0�nK����]
��8����`eaM��?��w3:��?}�K�w�Ɩ�����CG�T�V/�1[q;L��i|�^:o��
��t�\lr�z��~�_}�G�����wPչ��``��x��835��Q�3@��d�w�����:�x*Gg�?~�i^|�i^�aY�
���$�)�V��!i���jR�B6F�~��{�0���Jt��>9�ʹ���:u��-	��@ ,�`�<6���l���g�	0N� IH2
Hu+t�\U]Օ��9���zw����?��<�Tw�9����;߷���w-3��. ��0��ϜUzҺ��9�T�x25� 1�+��YaSY�s�U�.1*���R�U�&�]�f�\�E�P25_��#sI�KM�$c���*._<�܈H$(�zV�5�L��*T��i����[GN`��������7��E-F�^�ĭ���,�>�>t�.��u�'p��xcQh�0V�y�e��6،Ԛ�n�@�#�`��զ��Ҷ�bs�����!\��`����=6()0�Ξ���g0��G9O�9�|������C7���@��D��AOG�V[;XJR0��8�>,N���I�:j�,len��bCU�Dۆ01W��7�ê�P�Uq�ʤ$Vt��b%�NYj�xyp�(�I2��(��l�D��M�Z��SX,�i\������n��@OPN �,h�D��	�|�b./㎍%_d�������[
dI�I8����=χ�;s�0��}��cIcmvnx�t�?g�K~�+�W�t�<}Z�e��m�Y�p�D�O\����d�|/�V���*n<y����TȘ*VM6Z>�7���ˊ��c����1?s�m>�6?v�����Lp���8q�54������vI0��|ENjwә8zz:�+e`UP�����/ʵ4�A|���T9Z�&��aa�S�	��g1=1��Lq#��Z�C>�@2S��Ղ^+��P+�@)]Ɩ�8�Ҵ��ˋil�v+n�{7:{6 �� �*`hx�\�B>���ԫY\�x'�?�R~���0�2X]�q�=?�]{�E!S� �/@sZ�5k�qy�d|�����'q����Z3�yw;��
u�+F����iG�^��^��
�����i����b`%�E�T��*p�-������ V�\�^�$�
�a�Ɓ�����"�_YoB��Q(�1}m��=�l(����}�!�&�^)HIۢ2/R�m���Z:TZ2եt\j�H�(Ԭ��̓��,�̢TX���j��}.X��'�Ѱda�}���=�y�C��y�#�v_/*�������ދ���;����C�a��t#���K�m�H�ʨ)����_���m�<��o��Z���E
���H���� �A�̤3�n���EmU�l�{F�051����1W�ph��Y�]���:��Vg�E��<G��x��I�8�8�kpvщ�{;%ļ��c��,j��g.����
;�D	Z�lڼQ��f�4Y|��ؼy���o�YM!���4�?Ѓ\9��E��,����RQYB�����)��]��|!W�F���!���s/#[���b�g\�蜐k�&�Tje�Hēh*-tvva�{Aw�U9v{�l��+h6,P�J^��\Z2_i9Cv��d��.���u�n����Z� Yf�7]�#F�� �e"��ۋ�|�r�w�n�0�GSb�E6W�����Z����s���h���p!a9y=����x1�% ���2�|�j����ܴ]�A4�ʥ44kG����T]=}F!_���|R�f��K�}�N����췋泑�C-�B����;rY�q�7��cr*�ba CC�P,L���h��R�L��    IDAT��SO`f5�����0z�F����W�<�fA{S����l��;~������II�`cO�fF1��"r�:6��8��zK'�
��R��q�VP�v��|�f�X'�zO�x�;�g�"���U5i����J��/ ZB��Md���uCh���n0[�����X^�4��x���H�G� Hf̲�O�DƐ���Z�1�H37܈��lt�懀� ~xè��������
8dno_���u��2�ò/?�/b�$�9i4�w�\�=9�	��R�́�ܐ�:q8�0CM���^7����)�w��E�����?~��-%�jeSW_�����1�D�b�'~���=4X�, ���կ���cH�aUh�_GO��u&�t��{����ˣH��`!oL�2_Ȇ�#S���w!��aq!��Ş�7a�݀�X]��X<w�׮�Z2��竘�����ֆ��8�2��*z�=����R�᭝E�D�V��ǭ�=��FW����S�@T.�|첷05yǏ��Lf
����	v��F�w�w��jM;�U��F�
�P�qS�[09s?z���-����P�7�QmXNeEЪ�SX�22m��6��&����E\"�G�j	^���	��Y��v�v�p��&���Xɢ��'��V+�|�0�%��+2����q�2�	6p2�����1�l/g��l5L�%Au�@Cs W&�َ�H��͵�����5L�j�U�h�s!Yh��������g�����6����	
��^<����ʓ�9ݐ�YK��"�u�� &��a�v�:&&�P+9$��Cz�8�o�#�:��̓��[�y��L���\�0=���E����;��R�jqCs:�uY�K��[e�NK��%�c)UBl�^��v��v�t�7��F�#7���j���nX�|��#��Z���G������-���_�<�/O���λnGgg?z�Yl�<�?��������'�~�*��t��+�gԡ����N���������yly̌���s���]&S06Άz��@"�ƌa{"p؜1��f�\���u�;1uMG��AC��).���.l�T�`�\��^D��â\���ٛ��NX~_@Jhق�괷Ӏ���ZdYN6=��E�G�I0A�� g��z�'�#28�N�ɮVQ근~����,W�vt���Դ���U,P[نёA�{�-�?���(�(��,��)�uD�?�)&ǝ흸p�4���<^?[ss�X���-��n�eH���Hf4��x/}�����B2UBw�n<x<��PZ���������)���8���pX��t�mT�)8�*��`�zQ(5��$�ՍD���)\?��M�X���e���-�W��!4<��s/�X���]�j�R�,w��ł���Cд8�)p���x���`mٰ��*v=4�e����3�rm	��=M��{�km�oU��lܐ��eT��`�ϑ�k]�c�����pP�g��� �b)+㢷�G ���s��-���������$Ȓ��V�V�Mg���=�@:tH�,òD}��a<��c2~Μ9#c�`� �?�3��<7v0􉶑2��7�sX.�y����:�^2ޮ�=�Dj5����>XWǧ�O������:q���hf�b����$#�����O�<98�	���=�����շ���$�+6�D��XYM�~��3&������ل�/���4G��Í�X?�i��9%���ei<�O�`��!i��[ø�d�j����hY](���B1W�_¦�a�$PI�->%#�����w�{~V[���Ns�0Y%�E1���ba�WOaa�<�f��ꨉ�M	��-��{?o���#��z��j���+ ��˩y�����[��cK���u8���Pd��Ig��x�4��)�(-�1j�4%wE�����:�*7	�je���I
�s�!c�]��6�[����nVB�m4�b��ͅU���-���=�2�9���Nv~��16,
��&*�T���Cv�Q�$�h�׀t����`%�C��������l�~篿�^'"z�e��}�������r��}^�";�bN�����wo��߆r�@ըA18ytz��m�]��/��Rq�+U�Sv�I�\�Z@�\�R��r����-��
��Y`Q�T�F���X^B��o:�h-�a�PV�-/J�����g���>����?�26�÷��}��yY���a@u��y1���Gy|��x���L͑?��}�q|�+_�o���p�]��w߁������*��<|!���˿��:۰il+�7�����^/�{o��M(j�c7���Fa~����q�XN$q��T���wP���b1��꒝�I!�,�h��v�������J?��\��r`h�v��tU=����v�f��N=_A�a�� "Ѡ4T�q�dS��	
U������n)�Q������>�~��>'8G.�\���{a��:�K��e=N��d)����u[�
D��q��b(ưdM�N�u�[�a���.\�{JOKNޡ�(Jz� ��[p��E��LT.��R��"�YF��B4B%_}*;=)
/��K��%���B�ڀ���6�m^T�V���ظ�n�O\�+?|��tB}'q��Z)��Ũ��D{g7*�l��@eT��^�����ׁlb�F��z�{a�cd�(fOC�."0`i�v;P*��|��B87����pqnNO3Wf�̿�n+��h��N���D�g���dl	��d�(ضm�X���	a��A���m]$�$�&��4#�d��Q���d�E�P��f���!��惎 �?==}�eWz6����Xۢ�d�
A �&���ÿW,��a�		$)� Sȯ'N	CJ;�}��o��v���[	��y����<.?;�
�	D�#P�>�T#C�m�V���D��O^ R�㎽��-\��b%���D!hTJ�:6�tr���s�b��
LӰ�Ϧ��
�*�%��FiS\�=��с���T,�\�'hC�`?2�
��(J�2�n��D''f�t`5�B�����3X\I��D�ٍ%�� U��>RuXP)��4]���\i��{q��2"'旱q��{�G���a5^��I#�
�ۻ�8����ax=<�ݿ�G�~����ͣ/�j�`�n�/>�询԰�Ro�y�e����JUX�U<��?�đ'ഥ�{��!+����UvJ��#F>����4>�jb�eU���ҨV��&��4a������h��LU,�$�Q�d��Q��j��Q��.�|�8vx,~6�k&�#�������zW�h�����F�ڌV���K���3n����<GCXN�풰�W��n�����x����������w�ًFVՎJՃ�U��.�:���y��Hah� ^|�UtGG�p��q�uY��N�@�K	(M=��h�:�2����I����� ;\h�kXY^��:����l2��h�ԡZ��7ևټ]��aی�������wލ��n���%�>q���'P�[��A��/�~�3������_���%B�c�=��>�1l�>�o܋���g���~�����������6<��O �9*1y�ӗ^ÿ�˗a������C�`�K8��s(�. ��*��T>��>��V�U��A�J-`�X7���4�5t�A��yXmV�i���P.�OP�~d�u��wv��2�uf�z�,�2h1���.4��	�˨Ը+�!	�ުXʉ�@�X��۵��fM/;M@�	�.��7DjY���١g&���ߜ�I�M0F�!�lz�L�H��K��L��qc	'��aߎ-����չK�{�ZBgw�XD?J�:jz.'��M1���%�|^TJy�įax�W '�����44�4��V�.	4�4(VMkU��z10�w|�W�JV�~��'�"]b�3�pU,MO���T�*�#�Z��ta�j�ع�)h�J�o��D3��z�D1�ŕ�`f�8Bކd��� fzx^�/��m�JA�a�-d�Y.����U'�ф7�T���^�*&�"�!P����������<�v�s�*�J:�[-���Fͣ��A��c�?�wiH�Zq��1c�7����C�.����.elH:�}��4>�X��i���Ëj�&Z��ff,��躔�7�������A^��KƐ�����6�cww��]>��a�
Sv�=�l�s'�����ׅ\� ���U�Y+b��aX��z��8}
;��1J-���N�~q�Ί΍W�m��YM`#�GV(Q��g�`�:\��P2[5�:�����V�� It�x���P��!��a��*dW���X\M`f%�|���	ju���ۑ�P�&`5tXaA�@.�ò;f�]��~2IIC,<����0b�a�ʆl��TfRy}~�*e8lq~x����fO�"���b��\7��~�7QiZ���g��h�m��~f��2~��w0w�0"n�:���X��`eyQ��a��zl�h�o �<+�Hd�]�.l��Y���>`k��m����hӔ�pR��)����:�}��i棞� ��2���Je�c�}2��c��2;�y�"oh���JPH��2��)�(-�ΨQ�7����;�����^/(x�u����u�Bj
�O��w����zB> ����P�#��م+W��u ��Co��m!��vcq�4��E��E���.�|>�*�h�NCA�\E��߀͒î���p�31!0��ŰBiR��y�,���ܠ���F����Y��_~E|oz��$�(>��J��;�����;�+�_�>��_��];���^~�U|�����G>�/��<��W_��=�_����t��C��s?����!pঃ7�%�zzvJ���Y�m��n�z���^|ӳ?A���h�'R������1}u#ۡ���N��CGo/�����W^��'&��j�������C0 7bm���"O�\  ���~��.N�,�,�Q�G�$˹ܙ�M��T1f���No�0�����p������!�X�:�� '?N�f�X�Ԡ���ɝ2��1~�������mu��)�w��"!$VW�g�6t��|���b�5�la��=س������u`5>�^|�Y�)h��� 3�{��H��Ų%�/!�ށT2'��#��h��b�Ii��*H�&�� �k ��sPma��i\�|�����,bN�ΟC��D��o���P>YPaX�B9����-v2����Í���gQwƠy=x��o�ן���B������t>����'.,��zÉ���u��,6������#,�ݪ�5&�FfO�L\3��8��4w������Mٰ\����g��u`E�� �!�H��,;:L	/~n�u�d����Yy�!�`<��r,�H2��<20⛘͊E#�ty,sklra#T[ۚ������|9�8�p�����^�;�0 �B24|�Q	�!�?#�F��t�N�~Ь������{�N���1֩`�XF�B�D�(��<�5�?w	V(P-�n�00�F���oM�v6�&�G�-�	ƛz�j>g �U�a�Ӌj��tv�A�ed��v�VӀݍL���bC8��UBݷa�ԁ��C�,�b�&�°��i�*����d�@ĕ��з�����x�������@��E{�1M}*��6?&.�SO�#2�I��5���r�]��|�͇��L����1MJ���W��ر�J�Fԥc$�D��5��7(z�j%�m�t`8<�A�jqZ�Y�P���u�ǟKY��d���Z�|_O�!c�����Ƃ����ۜ�L7LW��KX@n.U�IA�ڸ�7Ph���G�M� ����yLðH���P� ���f�<;�B ��c{���{7��?6���w]�0�y:p��<n5��m�iI��5�H�(�bذ�V�O0a�\o�9���A�N_C|ao��
����˃r� �O�L��¥jU��Y8�"��<h8�sip;4�%Pb4�p��+�Vc�f%[,$�h�x၃0[��������s�l��6�;7��K�4����Ds��? h���_���s��u��^�_����US�;���|���������o�K���`綝XI�E�0��~����cX^Jbyz[]س��[E�c��>�[X��o>�7��'��:���д0��0
+�n�+�Yd�E�ڹ���N;�
�M�{040 ���)��ӊ��C��I�V,B��J�J�H �3�Ec>م�&�H(�����E��VN@��U�HY��%�u�"�(�X,ɢJ�9>��Bƍ���BO��C��xsr�$N8N��d�)4_gj�Tr9��,ބd9s�⤁7݈][v`qf���c~�VS01}����D�s�ݸa�A��y����̰vbזm(�z�$ҩk��`~y�����a�Z�#�a� �N���jAo��t�P���S��q�m����Ǐ��
ʭ��I��Nh�:ʹ8�&��w!�F���R]�N��I�FO5}�� ��>!����vbd�.�m��rN�Ͻ�pćj��- ��J�P/.].cx� 4}6-�d���_E��s�#&����tB�佢d�,�jk�5e�~�% ���*2�����e\�s@���M0�^�{ㆃc�@�@��e�Ђ�0�w� �j���A��G�0��Z�P"�XgT8��ev��\�n�x�i!c�㐑ܻ��N}�	zM0F`������i7����{�XrC�s�1�u[���B��n���!3u��q�C��@+�����Z]N�*����d�+(���eKbץ����j���H3W%i8ঁv3j���|JMr�[�͖�愝=]�T�%��l+�6�؁TN��tQ����P�8���f񖪲YҋE��BP�"$PX}���*@SjH&Rް���P��uX4�U]2�>Ь��P�Z��s�|��\nF��lh8�������JS�G>�BKg'1��/��ȑg09�
�J7�b�3���WP|1IAɤf0��߮�����f�-��U�	���vc��1�<~֐����d��>�v-��٠��d�IB01�,���5��ej�M@��&������Q���p�en��+�T��M�]��u,�k��+P�.�8����Q�oϗ7o~�xݨ������
���<q�[�ە�{��$��
Z��<�̸�?t#�J��ʅf&�`SU,�N�-�ތ#�^@o8�łZ����!��a�9����9�*I�8B>��{ᰪ�ݫW3����D�Z�C#o�u�D����% #0w��;�7���_�C�ڻ;n�NW�R�풆�ޡɃ}��x���W^E{4&��DrE�Eccc�fR(�X�[���{�Q�q!C��4�_�!b;6oۄ������q��),O����9���P.���'����`�d�F}V����*>��BEw�����Vg&�6�+Z�B��#�O�-Ҏh8&�l�p:Y��W_��o���^ei?��;�R�t�ٜTt���T1
��DC�8��M]��Zu�y�,�6�p�Ɉ%X`.�4ԫr�	.�� ��z�QJ�lb0"b1&��$�����,QrB^g	|�-�z�����-X͕`�&�ǵ��8�*͊��Bg�$�L�`�ZS�ɷn��5͇�>�:��?��hr�8�~7����x���+�V��f�/w�RN,j�oߋ�=�RYC���C����<�_�˪«�LbueF�W�p��B�J�xz��h0$́�M/����Zv�:a�AC�Ak�D����ٗ�\����^�ku���pzm��D�;�ɏ'OO!�i���^{�M8|.,&�ѻa�S3��,�i�{-�Ṃ D7���l�h	`"��g42]�i��8 �[g�ֳ���%H$�"P�q	=���J�,�+l$!�J��d���헿A�ɍ�    IDATL1�'_φ/�|uy��.cIC��w�u�P�^�*�^����73}M���	��d�!�{�����]���;�Ò��A��)�]C>�����c�=�Db}��������\>�cļڂnD|nl�yl��ͲaȂ��&vJ���#�ԡ�Ѳ�Qo���#B5��*�Y���1ñO�L���i�ؕ��6���	ۡZ[H�P4�5`��V��¨{q�ß��K\��pF�Pi .;P-���
�45���!�ƿ��s�*,�ؖ����]LM�%'�z�=O)�(�F��o��1)'W9������>4u+�z�����$3%RuhV��i�4�Ĉ:�M<������"�*b�@�aT�@2SD��?Z�ZF{XC�݂Ҭ���ӝ�φ0����-���&d}3��H�/e�湟�� �YFnz���lf9&�T�"��=�qM��-|�m\kx̧��8\��s�^�����]�d)���Q�﫪�A(v�]��}��q~����w_�����O'�qkc�^�RC��GC�Y6JXoAW�H%�����+?~�|
]���%ר��u��f��C����jJ��Ix
�۽0�)ص
\����cT�PUщh�
�*5s�@��G"wd5��)p��TRŶ?8Fq���x��S�;�=�ތ���+9�_���7b9N�TT�/��&�>w.�G4l7�Aʦ�4Y�S�s����H�,�T����羏��nuC���I�Ұ��W~���m�7��[ރjM�?|�/P*�F�����ڂ]b�]5���/��F�o�?��' �$M��2��8}�4��m���(F*���߆����q�W�k.���݅xb	�U9'��l,W�%�J�a#�C��a�.�r�����fI��a�R�E�v��̵�l3^N~���9���G��!�p�=���2�lX�c-��\����Z/IJԚ��o����&����#?�n�� 
�,^y�eD�^$��b��|��ѭ�����ӮJ��Co�!q9�X�;�g~�UX-I���%��xPbj��U5���%P3p�6�b�C���P�cE�"�5���y�	��9�T+�Y�,v�UCְ!�1�b����EtD�P�&J��~��*Z�ܾ�-�HJM`�RD��Df�-��נ�\XH�`�_ �YF��Djف{��8��7C����W��_��}t4��=(+3�5M���h��z��a����Cw�K������+㦅�qJ��{Wx��@��"�9�#E���K�&�64w��e>(!+��B��99~$~��[@���C0�qñ�����$/%=]R�f���w9��f����-1wk����7cɨ����I�i���A"��`L��R�<���������6�Ϯ"?�Co�#��qXjE�D�����]۵C�'��@G�v[�d:�u�(t{Ch4�r*��F;E1;��:��`�]'�I߻&,� �8�Z�(����������t��255�����%h�pvފ#/��0�j�bw��P����c��h�0N8~����}�KS�6	���E6��K�s��S'L ��:`�꘸r�?�Ru	n/e(�˩�h��x�	���t	�怟21�v![L��6���k/}�l�Q��r8%�<SӐ.R;� v���h<LZ"Xo�F�+�y�Ph&$��2���4����:�G��uPg6��2���;�C�_��6a���86��hI=��B�;�ac�؍��Aτ'VO֭��x$+�y�,,�.��n����?�������+���
���g����[����*��,�jWP�WF�;;��5��kp;8u�(��$��15u�QR�S�y� L��M+*�j�D�vdrK�%!�G�χ����	��%baj�4��uB麋�(�!��/�W�g��߀?h�7��k�_GW�l�.����ub˖�x�ɗ�uۍ�ï���8fg�L�wt!�։�>��ǟ�O|���M���Ћ�`vv�V��P;<n�|}����؂@��l��G�k�Èvn���С�0~�9ζФC΍R�����F��^$�e�<~h�!����v�r����m��)Jer(�l��G�����3��m�h)EQ̳�LxP��e񢫘l��Ф5��.�t�)hSe���!A�ŋ��YX��ļdӚ�1t%��B�e7}��a�xd��E#Ų_$�O��f��7�d����#�pmfJ��	u߾}ع};l���##�x��	4�yds	�/�K��ІM�{�R�af��sž�S��i���OA�$�s{;�gN���aU�s�E&mf-Kd���K����wm܌�N�uVV+ذ�4�=hٜ�Y�h���SX�����¦�� ��� �����Z+��Qɋ�����K����m�	�� ,���X^�{�*Ny	+�
�&:�7a����*U����7�}�W&�1>���g�b1���G193#����DS���������(�:P�s|<q����.��Y`~�����_\$��:�X��<q�\g٨`OK������i�7r�,�x�%���Ia	9Op�9����1�pr�(�E �4��� Y��K��k�a��� ��q{�����%����f�1K�fvѓ'8,KsA����*�.�6P*6��މ��^tvE�WSP��SGP(]�S5��,�(vdVҨܴo�zHgf�vRKV��N�'ZQ�`՘9Mՙ�}�$���4f�l��n���Ҽ�B���I+��海kVLN��Ď�!�wH����Qtv#=��	^��"g��Յx��������Q)a4J��O \x���矄/Dw�6�����v��Jk]�nK�:�N�ī?y��
�~����ex�Aܸ�v<��O�e�ðz���/P�!n j�"��N�|���O����^�H�n�_8|��p��Ȯ��4�WM���d�9�Q��HC"�Y�5BS;J��.r��+!�����[����6�Z�a7�d�����b>�?7�1M��2T�!�b��k��:E��A��}F��eB^�VE���hi�������]P��B�>����\
���������0Jh6 ��7,�e� �A����A��@�d������9ėq��p��h4Ӱڲ��vՁ�X;��3��w�J/]�A�����B�z��aפ�n��O��ͥ��_S����a�`Ƕ}�G��>y�(Ο��j(�V�BS��
XZY�/؎Zݎh�.�_�����%�;w?�������a����'p��Q���mp�5\=y�J�8MG(�D>�Ė�a���E��#_�E��­��(��[رrn	�G09q
��t	pD_��7,��F�]g��*6m�,A
���	S��`aq�B����Ԋ�:=~��>,./�PȈ�GS�̲`��J9/�����tk�,���n��J�j�Ҵ�z+e�ڵ�@G�:%v2���N�������䷼�$z��R"\N�dh$Q��F8���2�����M����be٘6+�KRz$@(j�q����!ൊϛMk�����4����DOo�� V�d������ N�~��O��ÁFm��bA&����k#�d6��,;�6�vv�'�WC˙�v��p�F�؍
Nc�LW�\D=o����Չ�nC�s�M�u�
�����E.���G�M\��q�m9���o�Rw�w`J$���e�/���,�s�[��� ��:ToK�����ر�vlڏRف�'���,��j�셳��g�uQL�]v�0p[��'d�֛/�xx��{�x�m]�ܱ"@�������Y�b��t�SZ�v�c�む���˘�f������l��g����#hk
�# s�i�d�M�������]P,��A4E���0??7|������H��l|�,G�o�Ɍ�&��=�!c����LAfҖu�j@{8�M���VRرu:��x���qe�(����@�;�e[�������l�ª����)`3�C��W	�lVH6qK�I	��eτ.�N�V�_������n��q��G߆�y?�f�`hd3.]m��ل�y72� �������*VGn�_X.͢��8�����"�]�oA[���_@*��h���`�~U���qk�ο}?z�%'��M���:������/`���Q�ƦPAwg�����_�+�x���af�r�	����[��+e��A��*Fr~S,uX�nB�Q�.vGF��[2#�򚚌˺xG� P6k4��$�D�0Y>n�Mf�u�%�u˚�:��3Mf� �%�4�>%븦i����Bi0aiYlk8&� .��BGRE�����X���.Sx=����Ș��ː��t��'/��U��X/pg�j���@��F��7�c;�+f�nO;N�:�
�J4gN���B�8�D|Z݂�ӎ.����!/��lHVu,K�pWl���4�T��"�����.ڕ�譪t�-,�Ѳqj<�_�����w��޿��G�G�(��=
�Z��<X�����[ĩSװ��G$lz��/\{.H^@|���V�F}8���X��wTC��ͪ�E_���[��`��10Ҏ��e�b���'>��ɫX�;�����k0=�������VS�CZ��+��s	�43���ۇ`��$�Z�������(�Ø�/��P���ǐ�$Q�f�|�V���H�W��১�GD����X�w�P����B�d�6��c2z�d\XC.Ό���	��Z�l����K ���fz^�xy�i��9���iKB���#��f��
�:�y�(>���q����tN�"q�4�f#7����hef�*��it��˂����pauuZ$�@��C|qY̜�zU&&�h�{ƶ�=�Eב�'�����K	to�w|���rG������k�7�Rb�4�m�naQ,��^jM����t�7��,"�ZE&���v�\�@��fq���������,�9t̟~'˅;~����,�AV�s�
8�sýȦ-x��9����%WL���a��b��%3�n�̟��s���?�=#x����{���{���a(-�O:�5M�;�+J1v��-�����{��wz��������p`@�1�-k|�����^;,`�Ԛ��:T6�Hgp��ñ��(��M4�v�fR7(<��yY��c�x�<O�=.���s�9����g�ZW�}��z�)��j�zЀ�B�bCw[;g/��?&����s��j��6��ώ�^B�\FO���(2��@UJ�f�sS6��qw9(��da��F�ՆS�Ca�j�d��M�ӌ�I�;̙��"]�!Ե}������8r�9̯�����{Gf�Ұ�*[E�+U�:�U�jm
l�i�=���!�k_�:�����}'������p��r�68�E@a:�����뇟E�0���!|�����1^��˸��{pσ����A�;�Ҩò<A!�@����,r�	,�]��[�����X8���%4�@���^���.5a�8?id	��� �@��_�4|4[�5:�u��ZY��Ϯ��tG�o�;��"p3��u�-&�� 4�#���,K����7�$84A!7��8��l@6F��w��@�j K�-Z:Y"�Fzw�黍&׃l�}��oPX)^��",�:-���*Q?�4�@�����Mغ�n8l�Ь<�����Oc�>,-]B�������@���׏�����X��k��d9E���,5��hz~ݘ
l�nc��K�"�(rH�5ܿ��ރ�ͷ��������Q).���ZMR�nԛ
&���k�mh��8ub'O^@�B�Ǐ24�n�Ks��_�4��.���SPe���u���kV�&%ʫn���3�t~�=�)�aى�~�)�yJ�{9u�|	٦�����"�j�.6�pP��a׫^��f�zA��K���Kn*n�OL�^���k))���:<<v2��d�����.�]�dlҙ�dsR�b�E8��!���o��.Yt���a��^o�ݜ�XTgN�	�k�ݻW��̲do�}N�`Yn�	6�(Tra�d��0??',��͛6b׮���zK�gQ�-�� |�LֈVn��d����'p���׉b-���6�jP*Mx��0Ҭ[�4�r�g��N�6,./c"uu���:�����\�zG^}��"�W���C���7���>��|IL�s����07���ea���P�ĥ���0sm
�5yӯ����s��%4K�P����}UkU�P��tL�W�a�F�ӌ���\507� ���˅z�.q�/��v2뾒uQ��ҍ�޳ ���x8����~���]�zU��&\��A'� ������%.�ҁ̺(��[������s��~������hq1ڍ����IsRw������s+������������W�?��Ǐ��$�x�Ʀ���:�+�'��0RR�FKt��J��.y��t�6M����N-!�cn�<�~7��C�AiU02ԍj%����l9��:;�铨I��Qh�&f���j�N0���ڄ��{P�MUϠ�Pmd-�Uk���vYeӗ\����-U��=�}�W����Kذ���`��
w�6�t~��J6�E��9�2��ik��r�~�5������4<�×��=�޾@qJǴ�i�N�+�q[1�p嗼���[��|�7���C�۷@�aA��@wo?R�K�mM�F�KE��ƛ�� ���λ�ܺw#���܅����^/��%%��HW0�y�mk<g�I�TAMg��)k`%�a b�N/�5��:��d������� 0�˦n���:(\�2^��	
�q/�*�A��vK�Vdz$��,���B�Y�4�n�-HU��)T]݈v���P��?{���
\S�y:��[O>^]�@�
�41��lN��XM�Е�F"ڈ���8�.��Td�ho�Bi5Ѫ�0�E�	���X�.:�J݊�L�
wE�GM(�?bBq>�v��v�P�7���p�{�~���'�7}8����alc/�6t��+�k�7b߁[1;�D �%f��G�ɉY\�6#�j�D�8#Ƴss�h��@ ��}ލ��ҧ0~�4��j��|���eD�A��{vݴ�O�����;D����O�&�� Z�8N~����*��
^9z��;0������]M"�
�ÃZ�$��SV��XX�B:�7���"���nH7X���bw�B�Z3�`�+����B�P�r
�MF�I�ґ9dB�bi�P*��E��QFb�Tٽ�����ǵ��4��62�dV֙����'��*�;��J���9�Gf SKh�Waa
y��qE�v"�y�ؾc#t=�ï?���0)JSEO��v˝��k�z�H�Q�/���A��Q��߉|1�H(�|6��@��NM !A���~�� =����AWZ8����ހ�ًM��ņ����_�Sх�l،XW/:{�$E���^B�TD�� �vɵ�����{�=��r��q�u�1�pY@����b>���@o���&N��ݛb�T&�H�XL-�Z��F�mC�fG"UC��b�ʵw�s��K�"���׷nCCP���^�'����+}%�m]���I�"�:���[6I	��h�BF'�t�,˟�8�*d�?`v��R�.cϞ=��>=5%���S,V�<5��F�20�M��H��2�
�|`1��c�3K��Է�������-�ؕ�{��~�ڬ���M@�N$H�/:��1yuV;u��X!{����][�q��T��q�-y��V�+y*�x��[�I'఻Q.Ђ�)�f���4�;�R�,�2h�%��6)i�v,�. ��������D:gACeb��r	A·F��,"�^�yj�`���_�+���#/��3��| 6Ja�nD5o�����l�o��3L���]U�v�\�U]������圈�LN�lc����c_8��c����m&H $@!����M왞�霻r�����.������MwUu�޻����� FT���Cn�"&��4´�    IDAT���,%�ҋ���v#���lqɨY�. S�0?+��������ȗ֐N-bxt3�p?��Ocz�<�;���M��:�TZ6Íc�Z.�N�	K���8ɉ�}�cl�F��/��{>7���H�8	�&��cDG�:9�m*�թ���� {C�é����N ��G����m8Y��M��N��;��z��
[Ndae����:x��[���t�7�hr�2VGFȬ�k�Q��Q�7QUU4���_�%w�uUSx�������?�{��Ja�v��ɞ�9�����ܸ���L��E�ve��*Ȧch�X�� ����-y���t}P�4�I��{`UMh�/5���,�P1�`�[�W�(��׫ x&����5i&�������r���=0�z��/��K����l���:.�Oa��kp׽Z͝�����>�яK��>�!	�6���׿���.<�ȏ��?>���>|᏿�}{�cr�a���x���:m���?/ ��sä���/�����/p�{;6@%������Oc�.,�M����������8:��Bغ�0ڃ����b�S(&s� u�t"��ceu��!i�XXLbj� ��6���+��	v`4�Q,f����]���"َV��\A:�:i�`��>��|^B�����_�r����Z��0Z+���!  h9�ؒi!�H0D�@Ƈbk��ۭ�N�)�����׊<��qzr�
�̈́M�G�C�w�"�cey]�.�>p��0ؿ�l6�#�[�Ï>���v�.�	��O��' �Հr��kz�L�Ky4QFOw� P�]�*���2��"f�a��U�Z1<|����xzc'^���&��n��I���?�K�6*�|^�Ka��u6nځO������8~�(��_�D��S��gԳ3p���w�{1<��<�f.���^z:m��d#J4���҅>�D��Շp$#��O��O���ثj0bu-���a��k�c�ż-z�^@:�9��3������%`:p����5�M�������}�Vd��"QB@pW(j/+��9�ٳ����D�ڹs�ִ����0~a�@�|?lV��_��57��መ��|�_�p^���|l$��T"-�5Y$��-m"75'N���j�|2��Z:����&P�2�o���lz���O|�#�f�vD��u4�c8��O����r��Bz��rm�.�r�I����d��\��hΉ������浄�j�]L�R6YL(s���D�k�4B��f�/M���f�b5��.�oۏ�Ί㯝��=
����lAf]~�mQG"�ӠB��`ק�_Fv�2��f7�,Ξ�@&d���������T�6��\[6�"�cq�"��<
�0�Co�#=��g�¦�nF$����.�E_��Z��hb��*��*
�%d�e��#_Ʀ�N�O>gs��,l6֠j�6�x����R78�ա�P�=��An�e
��&���Ƴ�	h����x=�Pƻ�.��k��[�עY�vpP��O��Ӭ��S��f��ϚɎJ/1��(�`�MS��4��y�"W���Ӎ���u��4���?W���\(L�����U��w2���`n��0d�	-q��RP-��Jב�Rga��Iglv�^Ꝕ�	�����,��,�vU�ł� k׬�̢)��HZ�lZf�I�����1zC6���|�,g_�V��v�����N��Ο����'&�{��?x=�d#����s�__�s�8��/~_��/��>��n�	�ύ	����+�{�9���?�>�y��NN�����vnƾ{a��d4~�$�ο�Z��T�]{�g0�q/�,��ͯ�X���~'���>�r
��~x{wbb.��oN�w�C�x���>�mV,�/`l|L\�d7����<���ϯ��+�U��-�Sk ��	�Cؐ������+�h�sE)�B6;#G�He�YA�ϕ�9ђ��0 X��t��cg�;�4�������JB�>���b	���k�I���(*��K^$�FwW��1?�_?���!(�:z����gE�w��W��g��=�-���p�O���6���`�b>�hx3�o��+ �2���.,��H����e��rd����X&w{�+=A�z����s	\��&�}#7�g�fT�<��S���/h�]�T%x�n3et����u� ��`vi7����e�=��o�k�`Æ>��w��~���1�u��w갡ۅ�P@\�z���#�?(�(T�P�6�~�$��g_�/M=��Y�H�u�|>��C�#��^�s-����(��6��\�d׎�xCnA�Y��ؗ:S����\^�����=7��m2B]^\�������"򅮮��hEU%�LNd[���k����0�6	@y9�n$ڈ�~����(��㘘�!_������K�P����bp+�iF��JRHe�2���7��kH��ºy�'��/�gH#>;���v�5�u��cLv��%tVlm@.ʀ.���9�E��N_��ф��E)U���u��D���چ������j�:�Y������@�
X=�1���_�Ň�v�����;a�van-�l&�h6��́F��n����a(�zڽغi3M�}o<� �f�0�� ����n��rIF���*��R�b����x��7�01���n�-vq[��O5��RTP���!�ǩ��\�����k�ǝ7����A�������3Xݩ��cxj�M�ѣ�E�H'r�����\Ӽ�b�\�d�%�k]3(#^�szm��w+R���75��	
e��z�5�������(�GP�	4�(T�l�{)��
�#S�	����C_߼�}�^�s����������A-7sw��C����ݰ�0%]���q�z�,<5��㇩)	�l&�Ao �XX�&�	f�MvF��aRpX�s9�;%���J�բG�Q��X�цR�)�A����U3�^,���> ׆x���mx+�6�x�9x�~�ML�=؅޾!���t�����?�Q���chpN�:������'0?��o=� ��⏾�x߻ߋ�h*nɘ��ӏ������Ė��an�ƳϽ�v�#z(���Q��~?�=�0=~gN=���_��͈=�v�Q�.ۉm7�pt�Y�`n.&�v���f@:������\� G� ���ێz]�w��]<��PT��5��b�� j%��*]~���e.�4���8�69�t�Rƅ��v�msad����z;x���s������q�\|�E�V�@����RW���E;F HvFn��OZꛆ��A!����?~���؎�|�K"fש*�8zf��pl
��y���!l��
��D�Z���2��D�X�h� �8^y���0�m�C� ���꒛q,�b0 �Kal�JR��@3�@W��}"���Ә�����<	�ɉ@�~a=j��+�x��ų�q$Ve+L���չ�p�زs.�L��$;W���)�9Jh3EO�����7�_�c�_E��D�]���fF��Mpwވ�{Q�a0��������~�b	XlV��z�D��	�K#M+R�@���P���@\�z׻\	y>M����
�1d|�ƞ�dd��,ݱcG��=���
�mn��u,/��¨(zq�ӹ<yi��S���n�=$zW����0�* �*ff��\�Z��f��'�^��t0`���cYj_i�B�5֓�*�>��5Ǽ>�f��g�`4��!��q��)]��e#�Зk��l�<��n�	�SS�;*0�. �H_���v��D�ZB���lw!���.�׊�^l�~�ˇ�J,I���n��������y�lU#���;Fp���'�A�.^:�Źq�y��h���V5��
�Tj������%<�O_F!C&��g`��Q��\��GN1#�Hc��[p�S�h����A1�����O��o�K��7up���	��m^��$l��b����P7n���8}悄��T�X
�]�R�gPM2`׺b��(���l|�l��ذ� �}�MH�?���W�t ���`Qd:��V��W����,>h(s��k�f��=��s�H��3մQq�����Rƺ�c^���o�iDC��t�o7���rj-�h�-�F�C3a�e�;gx6��Q�Z=�1����t5�h�B���[޹�:��֫P�Ә���~�..>�t걇j������B���񢰆d�r�:T�k�g �zf ��8�e�2�5�E5}��\�\~o�dJ��<V����5��fRP��Q3�ŀ��+�2�jN*��ff����r6�F���ի�83�뮿��i\8}�]ؾs?����x�~���u�(>������)l��ǟ�kǎ`v�2�����|��z'B]������p��k���{pڇ��nqub�>�߾��r���ѿ�\�<�0èc/�q݁�P�8q��<���^��17�]O<>;���OEa7Y�ub��nx��X^\���'؅�~�/p���
ia20e_�jE��E1-:���h�9.vd����.�	�׳��� G�͎z��u�uM -&��)j�\D�[���J���SS)tuuJ�u8���&S�!�.�i��x��ܥU���B����E|�����]'>�K�h<�$�c�_��nA4�G?�Y�=r�b�8�V���k�ņ�N�w�`���Q��f�㓚��ܼMF3&�/c��݊:���ql�F��Oru/{ޏ������`��4T�e0*�H��R�k��Z$��!�R.X�6��wލSg��ؑ�h0$�����fn?�z������e�|�$\�[g���@���j;.�Q���q�5��[A��`avnW�����C����擣3�#�'J@ZYj�QqKH<�����s���9�_�]���&D����`p~~v]K���;Jz��e��r��٩.�t�RC����-���d�|��10���`�>�V� f7�7"�.�vU��$��k��r�-��;vL ���&��\^�۶�s�8�=~�D�yKа����M^^��\5�Q~�"#�t���(�V���,¦�హ1��:��](�U\8���3��6�`'_GC��ӕ`V�X�;�ZCW�E���F�ϋ�@�Bf�f�K��#�{�^�婳X^<S��C����نP{�[vcq)ЁG�*�μ�D���~��m�死0<�	�l�.M��'`�塔�0铨5K�����@�Pǯ�}I6vl�!�ע֤1���r����>\�t�4dA��aC��[߅o����J��l:��<��4��]η�ǍZ	�Sh֋p	�T|���]JK� �|��46nDt=gR�l�|*�B����(4k��W�&�VLF�ֳ�ψ9��9k�	�DCMwqC'��ِ��f��&؇L-��FqSg�Il��Ȣ(Ԙ��d�d�[�-��l4���Nӳ����*:d%���������߿�]�w+W�\=Wp����<����w�tR���~�\�z2�a��a�;?$UCɢ]�4�]i$b	�U��$�[x-���ΌR� �� ���*��&�[$���T�E�x���Q�*��z��F��%�u^t�����Շ7^�?����v���'1~���z�o�-�E�(�k�t���»�w�}�8��ki��?}O>̟�̧�/���R˸�k���}P�V}�>����P$��X���5�q��}�����5a���y��o�i28���Q�,������v8l!Dc5�RUT7�u�m�y\X]]��PE6�&��k �vބb��B��\���΅��G��f�\�cu5*�\W�Qm�f�ܤ��!���`���������jL/w��e�*[Ox�j��!�j�hA���J�[#�R--�cj��;"�<��9��Mt;�"���$�2ͼ��f9<������Y�8?���	��F���ɋ2���Z�l� ������>��(�W��c�D����*p�X�k����vaF���;�(��拸y�!�F$s��v��u=�O��G(�ƭ{���^<��S�Db�&�R5�˕��ET��T��Ї?��_~��K�<�AMcn�$,�
�NFvߌ�߀G��5	�vw�Ai���
G�Wr�zzp�L�����
(�x�(�ҁm2r�jA>�:�����-0ȿy�	������E͌ʥ�E��t�ZM�MxNG7�˙�J?�"r�E�8?{��>}R��"��㢛��L����5J�n��M0���aɦsZ�P$&��fU
�Po��x�!�ǿ5c
/��!�Z�26oތx<
��& UZ#({�C��6���x�ay��s��_��Q��5�*��j��l*����
\Af/�@�[��A�[��?�*t�^��O�/���m��n�a-�G���vl���e�F4*IX�*ҙ0LV�6�VIYi +��Tд�Q(�qm���Zb	�����c��q��1�ڀ�ߍ�-{��P�8����̉�P,�����R�
�����|��SX\���`l�͘�w݌;��t���#��e��㫢u���,1e�=�.�����1���x�����ٍ�sg>yK�����ko��bu#S�5��m��`I	�v��������g��Bj���#{��,:B~ 6�
5���U(�"L��_\��-4��d|W%y�1��7Mb�`���xB�π&�!	
UijQ�ԫe��T;ڋhԵ�z�wҁ�:��ZK�\�u�t�7�{�,�uj5���)�45#���1�Ҍ����Yt�E`t��,�����o���[uX��S�9W
�ɟ����j��{�ˣZ-�VՁҍB>,��QqI�2��a��8�z���N�	��U�#_H�Q��is!�Ѳ���3u�p�$)�����aJG[�Z~;2Cg�k)�ق	U�����ۅ'~�(&ǎJ�l��F��0�\>!;N��K*�<���~�㇠W���'2ؾm/z{�5��¨Ջ��رw���y�4F�P��G	mFl߱�Ί�r��������0��Z�/"�x��8f��������\�.d�u��s����\!�5$rdl�F���f��>uƦ�qu.�e��ې�6#"�ʺ$:K �������dJTA2 <O\ ɞhA�:k7*.�dL��Z����c	([ݱd|���g��r���RZf$ѭ�r��v��[�����fx6��ߕ�"�Ǽ!fSiB�5<+�%��u7
�NE����r�::�p{=���C�T���Mh"!#M�q5p��K�X�HF�
�/���*��>7�V3R�(,����dղ���0���	�������[[BGW'�<�D<#c���y��Y�GG�B_��t��P_n��V,�O�ҩ�8|h+.N�j��SA$����_�����=�rvj�/�`�P-�P(.��aqɋl�%����p�<�/=riM���.�r���|��B�o�T�\��A!�5��S[�vz�����11M@b���e9����ҁ����$E�@�OQc�MP�*r����K��2��H�ao�����ytvt�&8#�Bm*�L^�d�����4���'˘o=���G�m�>1g��C�"���yv�K0w6%��P0(?�����{\��aT�V�[(�Frq�jAƘ�z#�&((��sw��p�F�������k�{(%��;��t�;p��BriK�ch�a��5*�:�\b��r>w&���m��0"�,�x�?������(/Mcu�,:|�>t����zr	sS��ʄ���/�g��^��*T�u���tv`���{�m��MR��|��2�&�!��#UHbvq�7"�ȣQ�������z3�n�m�m�|���&W�Q����%�JY��xK�(R�
*
��M�U;�;<n�zGq��;�ӵ�D0}��D߀ג�D
���2=@뫰�5+��\1A5�PoVPk�P.v�&a��1i��l�    IDATq��o�����˓+,�LW3J7sC)����`2�����a���G�1_M��!(T��q�M��ͼ����l�h��3�l�ih}�6+�L2�F��@��õ����o��U|s�\��bP8��Ͼ[+]zg��x��8��Ŕ���9��r%'bp�n2v�l��j����F]�\���R�R+�g�$�x��J���(�PѨqת���z�",j�t
��E8m>,,�1��l�uz�F��O�ŧ�YzJ)��dr�@���,�
E�����و�_?���dre���P�I�<��HD�d*�����5}�it��H%�Y`w5�_C�ЈD4T�e�����G�f����?��6 �:���7��m �Z��Ը�@+F�")�AT��+�����Ga�5e�6Xݲ#-f
���^���V�X��Y�p`�8P��9x�~4U���6U_y�[�.�~dO���9EU�=p�oCm��]F���>��k�"NZ@��! ԘI-��,2ACO��ܰ�|X�kҘQ)� ���2���(�6##�����p��_cr��
ĳ�d����ص{/�J��V���q��itu`���8�m[���4=jp��t0��������<t������Ɏ��u���2&���q;�������8��øt��������>jM2�i���������\)���lN#*�2#�.'����z�<A#�}�� �wK��g�dd�N�4��]���-�J�����k��jny��Kx����茰�E�TQ(��p���ش�A,ǿ^��lf�=$P�9 ÷����ح�M2�\���69��m$��(��s��tR^�����H"�p(fY	���l��a�v��-���C�8{�� ~2��(��V�Q����u$�x�I�5�d+%H;GgO�\_	ONNK�b�\E�ZXU�c�?�"jLeZ~_���6�3�q�d�IfP��l����Ä�.�"����O��w�����"ObraG^}m�.�-&�|
�P�d�VWp��g1��G1�����b���c.--`�5�`t�!�JN�
.\:��^����J�|��,��F������)�{��Ѭ�q��1��q��M�%�1�c[LN2���!�nڍ�0μ~�0�00�feg��aw� �s��5Tt�w�����1��ϊ\��6�d���+��m����7^�Nibj��n���4��׃�ۋ�������m@�L�
ο�C���h��ᵛ�JӤ��7<^���$�9����`�sz�&���c?����$#'�����Ix55�����&���C��5�ip�Y�R�F�|�'�Ո�jْ�r�������żB��	9�n�_s���K�(GӼ�R7/�H�PV�(�(4��� ,�ݿ{�;���+W�w�\1(<��O�_�L�[mDe|�w�f�q顢V6�Z���ɸ�4��핞K~Hi�'��d�#��
ugF�2Y�������*�A�RBEi���tM���F��JCB�N:uF,���y�;p�;?,�o��,�|�G��u!����ִ@WS��5D�c�u��g3Ν_��iV��M����#�j� ����H�ÿ�[�ڌx��'aDvgIz=�n�v��O��3�M.-��U������ۻ��
�^�%z%����/a!A�nB,_A�b����G�߆��9t�Bp�MX[^T�T�}nџ�21L�&��4������A��6՛��$�$W������|�o:�.zs�i�xAآ�����-����q�~\qoj�-���:E92i�R����ڼ��=�j���<.y�����yvz}Czpͮ���x��I@���� �<::������L5`v��4:��hԋH%���ED ��*w.�\|e���Z��`Ķ�M0�tr�^Z��J<��s	��[�����b����	<��w�J����F�*lGK:����n\X�P���\���"��,F8�V-@�9~�:�y��B`h?�O�"�"�\���z�.z˪R@$c���/�P
��kG}9��g>�)X�&��%Sr-����:!�+�9�>22"�I��:��ƀ,0�@{@�d%��\�948"cY��. ���W*��1n9>�N��ԩ$�oC����^mp�`դ%n����4�q��C��Ut���Ay��kG��0zIki��	�&g��j�N�QB}������Z�ߎ���	G4�jp�!��K'�Z,��cy�`4(���u������� ��ˈ�?���7��v�gx��E�H�3X\X�����s8t�m��0�L1�J.����]F�n�A���ţ��1H ��n�r2�@?��8�疥V�c�_?�KTP@�oG3�
C9�r!��m�p�����9XPB�G��A��A����G&���T���(4\�Pi`uxPEM d��PFff�$w�`2#]��D�l�"O �v�j��>.D��݃D��bB��䆂D��d���6���4D�s����5a1�3��bF&����̥S0ח���ൕ%�'W,	���7�v��sĞ'Ȥ)͌D��%�|�	�y',&#���/ع����R!-F:�[��'d�1-����[�T(Fev}3��.�*�6)�ȢR*��q˘�T"�a���9�f]a��n����G-Ě@���:�"�<~.Ead�P�אc��AA��{/,���x����Uhs�\��"P(��3�}�V�����\���]nԅ\\��T���AQ��H(+A�j8*L �t&���ˍ�p��C��P��3����ש78~Σ��p؄143�F�&//�[��KNb�;0��>�����'�c�<����#_X�2_�T7 ����-�\V��m g�MK G3��B�=p{��j�Zd�ް���,�g��L���#d��mA8���V�ݵk�9������Oct�^�M�Ņ#Oa�SBww�q4�f<��	���7	J��6�fՆ{��>D�	X�h��w������_@:E��E��V�:�E��EMo���͆D�pt�`׫ׇB���#\Hy�����	��Ӯ��&s�!���#`��s�V��%�Û�k>N��u�(���(m�#7BaH5��L��"a��KE������#3D��:���N�M�bh�S���H���c�6����nF0Ѓ�;����㘸|:�H-�V�F��Ë�j�dh ��
�W�!�<��7���ž�{�K��4Yq��$��yԍ�W���;��ߖE�PZ�c?z���)�7�z���o����"�8�M�����Y���/��&�6�f��(#2,x׽��k��@teS'E�����D!��҄�ס�֐�`�܍���؂h�x��g�~&�A7��5�\��B��E�h��~N�R'�b}y��������L'%�epp@46���[^b�u�09���:�\��fp�ͦ%���a�	C�Dc)�K�Kr���E}���Y�U*��-�q�]�G@��|�Ԣj#m�6�.��1<�d%�>Ek�I#	��l��)��a7��ܤ����1
�,"_��/������w:a5����J	��n��w��wcj�eX
�Q˭���D��N�C����3����?��㘼<���o���0�8U�D%�̹��ᱣ�M��t��/M�p�|�8�]{l�v��'a1s���4���2:�=�k��X^��`�n}��$ܹ��K��<���u�7WŨ^Y��Z�J�N�	��D"���ju�8���R��MpCe�V��`�s��D<C�/ ���Z�$$���ꈦӘ'�*7зi&Ξ��636�`�(�g��׌��,�7K2}R�**M�d3����3�0����n��|��%��M�"�珜^�ZG�FÉcS��.��]���a�D�
����QJ��d>'��Z;+���=�ZkB1X�L��$�f�vw����I+�����P�8FU:��X��'���0iެ[LW����N�\��lV��dI�d*ET�x�f�3�4�w������UPx�����LSH���?}�R����/��7�02��L!o�M�����qm�)U�����>�7j~�Qt��㇂��J�&u�k+���	����tyRd�יPk����QA�R���S(mE9K�F� �|���	�'~���D����� ǮÃ[��԰���7�TQ���|+kq���˦��AK�^�Q��n�]�݊][7�ܛ���_D�G�V�Ѣ�v�L���x���x���x�'�����C&�����o�<6��ѷ��t�g�"0�{0�i7&�&�r���;��g�P�q'��P`���z�=܏��<��W^�C4Q1����2(�2�3�̰9�ة��� �7>�Ÿ�ƈ-g�����#�qDt;�7 �s% �X|�qJ��rK[�o#��:�=�Ǘ`�8��f�Z��Lwf�*NS.�dehصc�F�����U�av�Ξ;���Sػ� �=v��#:6:m�zqR�tn�,�n��4Y}尢\�#H6�42�2���6�
'2X͗�0ّ)Աq��8xۧ���/?���G$�f�����6m݂�h~/v�=,#���9��,�K3M>��Q�{���u%�=s�F��,�,x�_�W4J0"W�	���|��e7��}����z�-a�xY%h�ZQ 3��x��rKF���x||\6����	�������aUu|�pL��-.ˆ�_�|���[�m>���KKk�37o�*��i�:v�l	��8��j�*�q�F�,�6\,�ш��Y�8==��)���}�p@0Ǎ
�濹A�k�\F8��4�#��) ]����J�72d+�����b���!���j����v�A{Ї**/�A�9�� �$�tm��}�~��FW����ގ��ưm�lڹF��c��^�G-G�� #P�e#��#S(�¨�}[wK8���EW{�.���Ǳ[C�oC>��r1�WE�a�-�}��;Q�\B=�"�h|c��c�uU,/���`���/��T�ȖW��y`��cy.��/(ӗ�0��F�6١ƙ��ZB@=ef��ՏT6���I�O^@&�C�P���A�ׁ�=>�Q�����Tj�%���7��֋(7\���v��b��X�.�̌v�67MvƗj�Y�okb�R����&WNo�߹	~��7[��|�	v��m�(Mʛh4Yw���Jf%�wn!�lN�װeiC��G*�,�$B��.��pl�'
�����K�!���He�.�a��eS�{���H}���6�#���*�u�V�X������������#pEL����|'~�Z���F���{ �^��.�oeS��b��&5H�fh4ٔPG;L��k�"*�9�(�K0Y��<�# �j�^K��PQiX�+�����˩�ٯI	0�>�z��tƈޑ;p����q��	�������ߋ÷܎g��=�������z��^y���J��L6��#���F���ꦚH�
L����{ �{����R��|�-��G"��b����4��[��f��W?{�z> �����'ŏ��7h�͡��٠X08�1p�m��d�:,N.�����6�o��Uf�-���m��Ё��r�k�u�#W2�o����ճ�� ��@����������M��j=�\��	�%C�N��Ő�͛E>F��z�;o��>w�\D�H2��@�u	8ZA�|.lX��TJf6�%_�`�7?~�Y���cg�h�h�U�vFGG��o����)m�,�@Q�b����=-u�{��G��h�Z���eL�\¾kvK�U��5]G_|��h��A2{�N�U�1E�Wp�3P�R;)�/c9�ľ��Îk?�|��������� �� ��6ahd3r���$�����p7�����3G���&�t�cs�XY��-��BЯ�©�Q�q���)�w��?��C��tm���,G�`wx�Ɖ���0;;��uca1�H4�ӣuhK�4_*%�V��#�d˸�rs��~�.)2�d�� Μ9%��c塡�u��&�b:��n$�"��-�܄����5�b���k�;��\�C3Y�Zϵ�&�T(hL������2\n�h��Rk���G�.|��/^�-ƒ?�1<|=��(�7�[2���6V�#�5$�-��(�b���Ir�m5��`�K4^��Y����a7����F��<N���ֻߏ\͊�~�a�#˰��݈����lܵ�̈́ӧ߄ZΣ�XE_ЍZ1���
B�6��N�2h�`~%���0:��ڤ��2���	���r��E���T���;����{��֊(�bpz��E��I�D�6��P�ء��%��Y/Ag2��z\�6�LM�������8
�e1��{�]��hq�h�Ag�Z�@5��F����Db�6v�P���C��φ�K�!�[��j���A�Ts���B�Y���3���)�[;� ��#R49K�o��AM�N��:̕�(.L�b`�V�E�X[Hc�V:��-�'SWӨ��B0�BE��HF�����A�Vc(W��ti:�C��hz��ڠ�0p���d6����vV�u��Z��2� �H�op@"��Q�8:",!7lj![�o��)�����ͽ��ܸ�o��^)$���+��N=��Zi�f���=��H�t6"�A1C1�d�c2{�t��R3"H��,%K'�<{vk��]���;BH�5�*5E� ���q�d�dT�(��(7��)�����r���XX,b��`��{�3�p��9������O����O>�2��X���Ŧ�;�x�h��?�~\�xF:f��`A4��>N:�3�(�2���/���!O7�0����Ag���nD��큠��<��C8u�'2n�����&&�W~�0��9d��n��wh)'T{?��Ū�3�u���q"[���-�dPpy�"�*6o؁��N���nd2:����q�Wdw[�p؜X[^�����ި��fM�8-�F}{��)����6�XK/�J��b�b
��}=���_��Xm��X�j�4fRc��nY�Ӗq:�\�U-�zqa�L���k��t�H����,(��S a�7�zҙq�eE]�MFl��������s[8��� �u.�Z� ���j�I/z�W�0�ҎR���j@�FѸ����Ħ}�cq.��}��Pz��V�=7���Łn�?~�����bE���k�O�$1+w�w�������s?�@�^Gv5���Ul���������ab쨌�$j�"��<j�4l�V�L�x9(^�=��5,0Z\2�"!�*�F��c�	��Ƥi��<�<�<��<��~�#�\�h _�TDH/��f��縣#$�,_��Ç�Q�9>>�9�mNē	���`@~._����vw�c�wM��v�A�����
uJsΞ=�dS�^e�,6���n���uʱ0�x�5
����Ԍ\.���/5h��z�Ŝ�ד��V��YG8E���Ӫ�J����$�ܠ�c�n�����[���ߋ��+��^y��}jŦ�6�����Q�g�7�<u�*j��#Mf�^4��k9�8|/�XEΙ�PőW��^t����|XKK�6����A�*gd��p�q��K����D"�N�͞�=[�����<Q�Wt�M6�32}�T�#���ZH�3��@Ft�s����ܸ���%���rA�/<�=��?��P���sp�R/B1���]�"�r�<H���T�H2(�k(g���݋z%��v����k&UKUm`�d� z�JU'`.K̨S��u1RhN�M.P6�Q�N�o�B~~���A.�[ �^qcv6��C�L��7:鋶��G�&��~���$����Xs]�)F1�qI��p�w�d7�}���]5�����th����p�����}����hr�]��bP8u��W�S�RH_*dd���(�ЫF�
M��&X���@�҆���8��Ad�9U�ke��,.M�@���ӈ�祭��R��3~�aq#�*@՛��ؑ�D�������Ȕ:3��R�^,�Ѩ�����bߵ��ı���_<�~�0��q�세��*z��`���T��u��7�7^x�lݺY�=�E|�v$itt�cq�2z�B����"�    IDAT#���Ie��4��<�=��=���7�o`T��������7�r��[�� F6�BduO��[0W���šZ�<]��8�@C����]����X�"��qC��}w�Kr�
�2�����ۆ�~�!�~�M��������9ol+QLe;G�F�5�w��^4f�[C�:�ZK��H�"�r0k;rEV.��\�[Bi��j�#>�R� ��XUy������dԚ3�Qtww r�c�6�Ȉ9�����_�ۥb-��H,,��kߌ��^�#���7�N �C���Y��|��&,�ܦ��D�����Ҩ�*�����d:+�{���E�oFl�u3���1,-$����k���ƻ�gU�8�74�W���_<�8=AT�idiq�Z�f�n��>�O-��g�@_�����hw��p�;� ������Kscm����{��7�3�O�Pȷah�:x��S=x�W���x="�KH���+7'� �xK6�j �Ǝ�����[�n]-ωf$щ!�قdפ�`��j�GF=!�����`�ݾ}�}�j�l���D"�_���pڴpt��岦seص�m�+���M���q���Yr&�$x��c<Ii�h4�%���.f�fC�8N�岰�l�c��� $��k�x��R>��(���J,"z7���Z���^�F��(�'a�awt���F{������W~-�ꣽ���mܵ�kQ�(��&��Kp �]A<�$٭�..̢���L޾kP3qqr�O@ɓO?&2	�ET]�'P)D��ǧ?�I.�]Ǐ~��%�8U.f�}o3ZQ�&�GNX-�_���h�ƍ{p��]0��(�<����ї�|�f'&`3�����p� �������Ȍ&��-���7���"�����N��㵋��h"�V��k;?k�N�t�2�?_(��Ko{9߀��E*��I�|.)#}�.RèWib&��AzA�N�b5���f���G.C���^��� h�1L����<��p\K$5���1��~$S1� g�)(�h��PL:j���`J.����6�}�\�Ef3l�f��v<�7�jY�&n@y�3��V����sCC(�py�%����54t�F�_�s��'���Bj
��{����M��G��|��+3��m]���h��oC"nB��օ>[\3/��h(��[v����q��8���
*%M�rx�J����p#����d1h@��$�����Ub�u�9]��q����pw��_>�7^���ڃ�-��������غu6m܍f� ƕ�N�c?�1�}}}��g���j�F.MQ{.�>����'��ك��G�O�9�W_y�v3�Qk�������Dt��i���v��1��������l�
��*�M���0T�P.�a�<-��9|8C�$Rh��D�YS��f��i��h�������cj>�ۉ���:��D����t G-J��>6=h!�-W&A��F���j���L3�hP��Q���|��kq�% he۵z�[ن�[���VBY���M3���H�Z5�H��. bue���v�=w���g�$�y&�dV�+o����0 މ$HQHщ��[J��=퉔V��;]�m��Zy�jW��-:� A�3���������������nH�S�OMG0��jS��}�����c>�ՕED��|�%�0"�`4A_?5nd�H��M������2�[�#�?���ט��v���(� �Q����%$3}�"�s�G��5:�D��AÎ������B��/|�����E!���P|��ë�^�[�ބ��!	
c�������|.x���z�,�_x��GLm"�UXow����'�����G~�:2qAU`�L�`A�Қ�r5��}C����q�K��?�3n���W���|>�>�%�D ��~r	�k�E���%�=��|�c�R)>(P?5�9r�"PF׫��0���xEf]�9�#1�D���ǣb��:�9�t���Ծ�݋�n��%�@�$tpسg3�ss38z�(�'/��23�t�����4�����s��;h�6���Z,摈G��s�cF��6����.�l�G �t�z��j����)LLO��װ0w_����ر}�&V.�מE9��p8���C��·�~/��֗�pϱ��l��}�"}(�k��*�\$&��)ʙ4x/�]gqs.C�����xam��"�Q�^���:���Ш�w�1<�����~?y�e���0���H�bX_^�C�P&�@�٪3�n:��O�ܯ���a1��?��?`����w���e�bid�q��^�u:��-�ȕ7�ut�
�[�~����E��u���t��t��z&d%��h�6t��ӂ*l�v��_���v�5���4�h�k��Wh/�l��(Kn��P�E���Σ����t�P���ErRk{���ML�O�Ѓ�'�J���a������:2d�;XYV�M��f(z�]3d@G��^t!k�:�b�w��6��FM?������ku�HT��E�>�d�V���`"�h���{x��?�
��H����}�(���K���v��c
�R��u���AH�"���82tӏPh ����շ���݅�� d�p��;0���Y��
}^D2I�@a	˛�[4����]'*	�J�YC����я&����~���{�Ǹt�5�{��Hd�cn>�kWo������0׮ϰ�k��w���rdp�7�丼|���H8�O��8|����&&�M���}	�);v�
�uܸ~}	�s���'~��Gpk�,^}�)��eXv�d��a$R����j��Hd超�B�c�!>��~ܸqz���J��(��;)H�{~Q�'�=H�IZ��"R�8�����q���f��L��&/R�t&�v�H�b�10H��P��vS�)�����u��>/��zc�V�����:Ƈ16��C�݃���x�g�H* YC,�Զ�P� $%�w6�l�V[G�]e]�����6�OdQZ�GX�C���n!L�|H����R�5ē	��-"����>���O��[7q��!N���Qh"Nar�4�����?B?�gW1�F4�@�QF���'�8q�^{�u�;�;ҍ�<"�"v>���D �ċ?�*�n���t�wa|t
�s��݃�<���wA	��Y1�<��_���1�m�7BG�����V�$��^k˴Q ������e(��7r�'�-2~е!��Y6j*iy�qE��m��._��9��Xz�GMȪED�I
.����v����I�B�(�Z��H����kF2�~X��
�����A�f�"P��Ԥ�\���*O����P(5ܦ���ٵy$MF�@��	)�gaR���`m}���d,�?����P"�jyg��>R�U�[�m�8z�q 1�����Q-桸��}�\��'��s����V�׽Ǡ����e�R�h�tL��AǕV����V ��Mf���¬T"5�_�׿�yw_��?����m�1��LN1��e��5�I�l"�@��,���c�ԧ>����;�>�7μ�`p ��S��P���`K�71�x��A�@W/��N��O}�0���s��<��*�jy��?T$�$~
�v��4�(6YD�MI���Ƽ��*sEg*gV�������@�!J��� AY�" ^:��ݥ��bFβ\�~����HOH|�H��(��˖���S`kH�ڤ�$��5�uL&:Hl�w����MPH�c���]�B2����޴&v������͞$��BZ2	$2w����O�
�'PX������~�^��X0@�1�m�cR�� ��84e�z �OEK'���|i��@Z���S��؝��s�Q�.`߾w33'�iA�sEΪ��g�!���<�SG�!	�[z��.Q��O4;"2����� �^�ዸt�$����˯��D4�#�C��!����o����w��V.�M1��I��d�7�v���|�I|�g?�op�2Q�W��s�  QCB��q���K��P`6O2`}��/`��P��������1	����QF*��U�X�c�&׺e(���o��-�~�>?�z�T��Eη���JN�zQD*;�h,�?��Q�|��9\G��ԫy[aq��n�	{a�މ�>��k0�ƹ��Z�2q��cr�1���5r��!�XxS�F懭8�!�#J��e"�g3�j��w�ߩ\*AE��9��a\�t�]E��U�atb�Ap,�F:5�c�h,�-�hca���T"M�]/�/����lԐH%�!��?��M�s��V�$�^G0aG}��Ɓ;���`u��ן�.&F����H������k?��^�׃d	�P�P��5���<��8�<�|�y$c4?�C0���q졏bhx��`7������(�ʀ�Fݎ�ܬ��]�";�����������(󈦓���Q�c��"����$��k�e
�:�u�kAt}��Lc>ό��:�j�F�s5~,�e> ]o0���CҐ��o��:��]/����s����|����䥒Id2I������[�Y|�]� �[�np���֭[���l� �sT���{�Zi���ٴ�H$�P��8zV�J�/�A��7��bPH�jӲQ�T�70�F���"�p����_}�12:�KW/"�|c�<��Ƒ[�⎟y�������%t�M(�|H�d�5v�P,��9��.ҩ�
ηOE�h5aq�-eF!
B�$�ڐI��E4.�k���F(A�a���G���5\�x	�_�!��b������F��O�T�_��J�e��v'���eC2r�~�����~��kX�m�Ꮋއ���d�c�I�+�w��{?��7Q�߀��u;rw�x��Y�/?��ٷΠ�Xp�e`���g�R@��eW7(��G#\�c�H�H6C�*&��D��=��b!9d/�YlP�*�9>��(k���n�T�jNb	),�2p]@��O�fȴC2���"��}B&JߠF.Z��St���&/f"@=9��!�c;d�r?MfhR�������hB��s�R.BM$�RHfO����鶦��E�����A�3_z�R��p<��R�|#
OC�&�j&��Lq��zn�F�Kg�y	w=�{�xn�X�����%!�n^{q��1�x��o�uL��u���H�;�'���f�`1�bw�������MXn�~�G��p�� ���g0����|�;����1�?�V�ľ�Qo�q��;�c���)j���t��4��f�}�0"�8#Se���,��տ�H���~\�z���?���������J�<>��?Dvh?֊9|��EH,�1�Ŷ7�EȈ���ށ^3��N`prV�H���O�Pm���w�B,��\�@��F,5�����Ub)���9����)�J�E	��5��S����ŊN�[�P��(�<j$�5&$feK��O5�[��-�";^/8�Q�x҄z#>b@l��J�W$2��~�,O[��&#	�ݹ���������aj*ˍdB�ڶ�k��R�R���78�\Z��X
�������^�]���-�ȣ`i�{��9�����-���&�7�	"�6N<�����tik7.��;�hio����''��/��o~c�[W�(xc������;�o���_�e�a�ԫ��5����e?z_����<�z�:�n�MF��q;�@Q��+?|k��{v݁�/��^7��t����G!��(��8������kN[��_��tPX]]e&����X����w9\�\�M��:C�\�toQ����(g�ni���!�����B
T?t�G&�;w��uۦ�f�H8E�R-���̙3��@'O�d��5 tݸy��A�eR�*Ҩ�~Ƿ�>�l�03f
�v��G�ӂ_$Mb��ŕU6+���UְU�N"ȕ��-��fS�0?�c{�arj�ﷃ�Ӱr'�:ކhfbr���/|�y
�+��2�R�`hb���X_]CԯB�����(Tڈ&�tj��Q�
TDD��g�4Â#����%���~�Y�R�ſ���Cd`��A����HG��؃H,5�@�|�+��2_{�9~������m~�=x��w_�6���8tϽ�8I��ף�9c��5�s�X�=��g_��p��<���~3��	���nT��U�"(8�6�@��c��Nw��� P2��g�IB�����8d�)�s��Cױ���M�I�G:R�u��j�p1|�}�5p���EC�O������ҳ]����!�r%7e16K<ױ��!��	��O��� ���<�	�Xz�hzb��B�&C�����B?�T���5���`�	��O�Nj������q�O�ǿgPx�����z��C��;�\�Px7��8ju�;�!_]C�/��׮b~�
��%�޵{��aqaj0���y��1�������EH�gC�-��-���D�mT�EuK7=L����"͋aB�+�!%�?��_�_M��^��7_�2��v!38Ơp��Cؾm/��Ht�9Y�B,m����o\E��2�SY�b����g���q��X�y���dѰ�9[�^��,����{?����������_#&�:Э:\�IN���*������������f9�~���zԏ)��5w�n.B
N��!i�om�Qs�Odh8@͞~fK���ܦY�"���n�~��iP!�L����:X��#}����n� =���7�75Z�Q��E�ϽP@P,1�ԜAYq�Bm6�:�|ߣ�����C�X���N�5k�������\��dF�hcn���]�3`4��Y�`��3�T	]n[��(�V��c��k�5�
����'1��q�B~��gѨq��MX�;v`vmv�TY����`A�z1�u��k�/sˌ�w�5k�i=D�A��E�S���羈�^Gs���9h�	��c��*����E�e�+��!�H��Ǳ�Xî��P�a��-DR)�uT�u�"Q��Ґf�]~ �2fl=����K3�6y�L�?�iz<1��ȑΕ ���ʺ��q6��F�葻Ygu���
P���`?��J���h|L, 1��x��:QDW�<�l�Ξ=ˇT
�&W��+�6!�A+���Ev�yd~n�% �cu�Ѓ��X��'8<������P�o̰�4K�X�pCS D�Vg֞F�V����<��w�8�'���$;��Bj����N��\;�C�g�У�*# ˰�u�	���H�u�(�Յ�8}���`؛zH�$���0:=����	�CiĢC8~��1�s?v�������>�w��6�!�R�=�}3�s��|������@�u�����<�Xp���~ۏ�ŉ�?S�C�R�f�l��mth���\|��8����>�����p��gQ_|����
hm�B�]�ȭ�#I�G5��W�)��"����8���T��t��M �G|,��(�b"�f�F�>�&��{�E,�a�F猢A?��n:��PZWh��m��xnb�6�F�֦V�
D�,�鉌Xt��RA�<BϡOM�<�hq =�"h͡�y�b܈}�lE�]�T�У
R�DG *�Tz/����~+���?=r�WX���+��|�($Mṓ_��v�aʢ���``��=�D�r�Z�t��İ�v�d�!�v&�����~d�Y���b-�ȡ��|�Go`t0
�_A*�"����6��\	�+E�Z�G�Ó�B'�m��I�Do�ܓQ�C����}�I������3�ᐄ�""�4�]�R�O��ۙ�$g�=��^��D�e���u�z�e�ke[���Ɖ�\Ѩ�q�XX�ar|�2��9�B���3�+���{�Fim/|�K8<@O/�m7�H
��� :Bo������;��J~�`�'�p��U見];�c 1���z�����    IDAT��ܘ��̹k�|墷9�h��"�B\�:�S4���vZ܈�����m��l��[�d��<��^Fe�]�	7�l���c�@h�q҉�����H��S�cl�k� &��u�B�*���w~��!�D��p�fn]��3�����ؽw?�G��4n۠����-��6���� |8��WP/�b�O���$b	(����.5��}G�bgH�M7]G�� �����O@/4q㝗p����54�r�f�aP�#�K!��G�QEKo�FH����C�1�E4���.sU�݇p������j�b���h�o!1އ��%�.��}��Ђ#�����ɓ�m ��mkȯ��C��"���P�`�Eun�H��
;j���1�\��zߪ*��IkJמ�m�d����	�&��ˇ�F�5�Ġ����+سg�f3����k�j�2Ba���`^Z]cз�����cã4/��78!��5��
;���06N��v�ƛo�aP��)<~�8g*��yמ�����@"F[�s�M*acE��9��AE�`��E�><v�.�d�1���tf�����P���IO,���l4�=�qTJ0�����!���W��C����X_]����F�J��Y4�6�qkF��T<���E���j)D*^��LZrp�����8��X0�l(�Dt b��/��(._=���x#�p�࣐i���q���� ��*�f	~
��p��[8y�{�e��+��������bϝw���"5�j��7Ь����.A[�b����W~������c�W�yED�Uc���AqL�ne�*^��(0-��ĭ��*O}���ؙL�?���/IC@̆K�w2U��<���&��PO4�EJD2�)J�y��~2Q��[iݧMӱE�w�I����84�g0�t,S����ɠ��,zYmHzjZ;��N�&/��,�D��W�)�±hD��!�"A
9�ٳQ��D�n����=�?�����p���+��|�3(���מ2�s��.�u
?>�X���Cp��B�]��+�����	�d�\:�T�6�e\�x�v	������l�\��6�oo��ܝD�K�E<7��o�b���e!��i�N��K��&���������"�(l��羁t�Z�p��;��8.]��Wgx��X[�4r�]��=~1�n��Ęɜ�#ѷHݠ"4 f���C:�ᮣ������z	�/��B>��]���]�1;�T�z�$���Z���\�!:78��]��\���T�޽��6�Hb�kKX^+p��}�,f���!�(���;�{�GIӗ�gSun��c���x�1���Ď�&G�Y���k4���6�6��>�&��ʐX?�zUu�����s	�q;EG煘��"g�Q_/����c���E��N@"W,x��H��%m��c[3Rݓ@�T��+��,���0�&N��
	�n��`@��]��$��L��E�B��ؿwЕ�,.����T*�E�Bo8Aͫ��JF���)���,q�nʄ$k�4DR{����E���s8s�ZF�:eB��ɇ��$�|A%�(xI˖��p��ETH�%�p%e�c��;p����U���қOn�sKx��<F����T19u'D1�g�<����apd;
�6�][C��F�P���*BQ��>t�n�0cHב��:��߿�??�4EŞ={x�Lן6�|�����"���=B�C:Dе����ueɸE��T:���K+XXXB&������{�w��p��z�&����w3�G�<
�~��T�U�$�Ţ<y(��J:��Q�wk�$Yf�KLjwy뭷p��㜍�j�0П��������B�ջ��/�v]j@��sVd֘ʁ�sk%���P���v@�u\>�,V�n���8��y/��Y�WV�IJz�P-�#����ʌ��s�r�2��Vk�*�����Ji>�n��
߫��)L�?��ڵ0�z����KR6��q���V�8����.��{J�F���FF���-B�Y<B���R��^{�j�C�8���ɗ���	y�	H��(�,�
̖���4m	�Ө��\��W��sw�߁���/��x��g��E���j���HOj2��$�|�d�w�!�1EG��Є	����Z�X�At����#(�+ܭM���q�>ْ�'�s�lk�F��Z������ ePh�f%i=����!�lt,��vz�	�&��0t2y�-���Z��%����|%6�ֵ-C
Oal
�s~!�Rʆ�g6��:
%zw`��w�#���vx�?	�~����{�߉-^��S����cu�4��܁x� �\GA~���l�It�&�\ywۋVe��'�v	#C}�X]@<���4���f�_�����et�K���U� �H�I����s��(�;TuG�IF��B��!�C��/}���z��hBy�>�Ǜ�_�q��7���e��3�R8v��i�c�����v���a�H	+�w�p�@=�����j1�d�۶cc� MI"�̢�,1�D��m�W����/#���;M�.Lˏ�k.��4���,o4�p��,��12{u�B	�M�8vm?�D4ź&?�%��������F1==��69CM��J0SH��̄����*5APO���b^_��	��F�:�i��Av{��l������h�'���A'�Fmt(T\Q9b�V���S��d��'Rk@���8D����!��ŜX�Z��zū�����29���1��k�t�4԰�r}2u�O�o�Z ����"�{��0t��ԯ�ߣP�s�QX;��SY4�e��M�� T#G��QX�(�`wKPCat�$�H!=v7��(��q�t�4�!�H�%�w�؏={�`� }/J���/���k�]%�����8�x6�y���Mq$hq�����1�W1<��.`c���~���,��o�F�}��J��_��� t%>r'��2�]�b�_i#�����/,�(���ڑlB�z9��q5�Z�Y
r1��[|O�m5/WM�v��G"�d֗�tM	H�G�bI�H�4��H��Xș[s���q��f���A�##ԯ�B��q/u��S)"a���"�0�
�C�gZk���Qry�*9���D� ��L?x(��#� ����ُ�8kq7�4/�B���/a��I���l��zi��p��sX�u��J��ӓ�:d~-[@�c���k<�ȑf���$�?FR�!S�^<��m��9h���m#q����'�ji�kd�	�T-"O��v�i)ؾ�2������?����}�	vY�h�]�k�˘��Hjn�7V���Whr�c� ��~��#|�$������:��TC�F�Ӯ%�GT��.5�\�!
���~�!�������Sȿ�5�����G�� ��I6Ъ6�H�V�4��#my��ب꒓�"B�4���z��Wf�|�1H��hB�-;=��=Ns0�1)�=Ū�pK78Q��H�B��=>�$%t��ѣ.�[�M��G&6��E����'"O��[߫����A�l�#�o�lCo��c�k�����I��py|,Ch�awp����c��6(�����+�A�ҕ�}�l/=J������c{Qi�+���i�7J�%ھc/��Ξy��o>�zq_��?�`5џ�JmG��h*�\N���6�FPn`xp�sK<>�d�h ��çFQ�6ydTkVO��E�+ p�8v�>58	-��
oD�m@�St��#S��6��j#����p��J�j��P8
�� A7��5C���B�!�cph�F���͎�kKK���Co�OJhϞ���E��%Ȓ���"�!ZAl4d�����[Ŏ�Q�ePj��<�M��
��h��ع}d��|a�5A����O!Oaz�4����^p�R�3�$�E�V忉@̉ɣ8M�T��ŋ�)�f|J��ch�:g�Ee�Sk5�  G���J~���'u��	�~OD�=�ml��^7(��}����;�;�&V�Q+�cZ�?�~���>��g�7Z*lॗ��Ra>�@��G*=��z�3�޾�U|�+�ё!|����y�:��g �[F��C"�	�I�Ë��cRQfe������m@��Q�%@�G��`qy	�>ǎF"����be�z��i��u(����C4Hj���,Q2{R�Μy�d�C}�|r���ݨ���B����A#�8 �+�Փ�102����߀����>����1��Z��8~�*��D�(���Z��P��l:�@د�A�ޣ�x�+��g���Wu=:H��v��=��P�s�Y@�b��F����������	��Lϡ14��
�;~�!&�����gp�=��H��z��ɤ�_Y�^`:��ʤ���aw�PIk���kx�YsH�с�,VV�c�X�����5
�q����6ܚ���2q~fP��(ߢh]�f�?�(�t�|�E4)U�~�SGV#y�-$bl�;0Օ�Q�";<��o\��j�B��A ��l5�Dd��U�HM����m�ݬ#ؓ�MePjT�8����F�P j�X%?�:V��/9�~�~��g�j ��*�<�lEbG/_�������l��h��?���?�5����������Sv၏�^Xi"����J�_�cZ�����d�B�]���`���{N��O<�N�&ĕ��*p�]4����c#���(7��`$��k3x��]ȊƚobX�Z�t ����J��|�(��]�Ůi���q85<�$�������&���)r����J��E�;�MH#iO��LUtrE�B��{���DN�`�r7G�4N��B��(����&PH� ��!���h�6Q3i/��@��~�w>���n���
�n?�=���k_�Q���H����������Rɼ�?���j�&����Lг�����Pɰ�v���D?��ݸ�@`�#WZ�:�)?�� ���\�A�M`=��`�X8t$~ө�%A��B��B���Y*�RP���f ���zOU	��C�Ӏ���UZ�p�bc�,��:},��s�:���UR���:$UC���i�*h^�h,@*B�T�O!gr��0�현m��j���ӡ&$��Z����X��9�U�"h>��X_. ���7`�4;$���5G�W}�Y�޽����W�E��U���X^j��&���;9��p�1�Q(1~ϰ�{�)U�mj�8R�u��x�
��)`´�G!��Z��F���n���kI����.z~/x�E���
j� ��l�K��L�ʤ�Ѡ�:�uB��v���9|�un5*��'?�{#!����=��\�}�����U�st������x4�d"£��ի�����$W�{�ƔV��Z&M��D�5i�p����Q�qǂ�`=H�3��<�K�ð�8u�'ܐ����j70:����(4EY�B��T �t�]��r0����%�!ܜ��k�peh1˗�����;1����\.4|��>�L����gq��"j�:�6A����T6�p$��F�G����)�kBѼ�01n0�ܪC-/�VC�(V<�!�A�4�%]�X,���]�v��fˈTo6�^�Ǔ>q}}�7H:0����=�-������>4�~��b	i��h��3�Ha}i��V58>��0S�4��á���r��~���m����7}J-���~W��$S�nx���XoL�}4�&����	4=��z��̱�7��1<�Ǌ��^z���6�p!�$tz^����id�qh~u��a�����o��Gi=��@4 �ۮ��q�?�xDEH�?��	��v��	��(��-h�.6r���|Q�+��9.��X�X��bb�>T�]tzn��k������tp�̏���~z���Q�]ka}�D(vw~�����z�aD{Q� v�9(ATm��!j�B���v.!la��0��~��
l�; �������F�͇'�nRЋm�.�F���F��u&�F2�����`$y���V��=����^��b�#�uh!��IZ��ז���mR'�,A$.9蹔Mh1K(�x���͠�&,DHzL$�ez��MPȆ�MP��i���3(�l:��s�	5��"��$���$��[�FJ<���f����{���ۚ���?(��n>Oư�na۞'1��>�u�R}CP}��RD���[38}��?�VuKsg��u�ba	�j9������4H�0Z��I�N��*��j��@M�@:��[-��F<�>�򣍹-���FG�1�&��%B��=*�9��z��Ԭ�|ڴm/J@��1�+,�Фv&���M��[Ө�k��F�jv��"D
�F�sxJ%�.TQ�]���	ر=-�C��GL	����ڶ��3"u�ҩ3�׏v�dϱ,t,�s�h#4[&��8b	bZUl�ְ���:Hb��R���>�����p
K�D�	�}�ݨ�j�~�o�]���u��KmH>/�~��)k�5�S�N�2��I��i	isC��ܸ�POt�c3���_�0Q��nUjl  E��J�yt�	
�A�)�%Uf&�T�sOq8���۰::��8&G�pp�6�u��.���9��N	��Q�?��Mt�Cxlr����f���b~�f���:�j1�ڞl�k+9�{t�z"mB�i�kR��ʠP���X�G����DP"Oard���Z"�6�@k�5��tJHe���i"ݗ�@_
v�	�cA4	�PQ�i&�h�t�KU�e4]ã#h�4��,P�^C;��K���UĢi�)�:5(d1?[@_���#�X��$V���nw�J$!�d���A��d����"�4)���T_�F�S :�6S�vd�9�b^�����	<���L�f�gUU�:˫W��G��|fw<��V��gt�sI��f���h"�d$������?}whd�j�(�PD:��&��b��CT�T�'��TB:G�l����[a�tPQ9ػ����F��l�Qb;�X0���,��P�*�������5�.�l8�"���xpp�C�����硑��/�Z�#x���q��I�����(�.$�8�m�5ĩǎ �G 5���N �8�Z]�G�#p.��	5 ���E̬����3X^�l�	t{��V'�����F4��j! �n��\�<������&�Z|b
}Sw}�IT��:2�AO�ҬqHt���@g�+�:�������`�:ڒ��B�	�*�)��4t���SC ���X0L�E��ѯ��adh�Gݔ�'����"��4��宒DE�@�5�n76��&�`��c�'*2�o֠ѡM9�i�FqD���������2�G�2�x�1��Fz6��od�{w�Lcb�^�Ǧ'z/��&T�����BK��d�d��o��?�
�+$����
i|ܨ�>�һ�I#� &�����G�PX�eZ��н��/�-4͇mヘ��6�o��*v �<���o��Z���P�0j�2���1t�9�<�t{��H��XʎU�\�#0 ��2}�ܘ@�9�]����l���F����,�i�E`tH���4_)B�l0��2ޜE�7}t�t�G [�#%z$����Z-��ep��7*%�P}.��5�q#J(�33��_�ٓ��ƕ[3��8zt/�U4�UԊu��Dk+���L���� �zZ�D��l�R�����x�^ŕ˘ڱ�v�;������ѢM��X�:�KPT�m���E�4��͎�P~��.��I{�;��Ґa��d?�����?:�BS���.B0-l�C*���j�:_�"�-�I�BZi�#�|=(�����4C:1b!��\U�`W/^������zu�X��'r�)�Wq�{��nq�OP�����i����,y�.��*��or�ÆZ�)ɵ����q]��&K��2�cQJ1���@�%�5B=�U4̅�}�    IDAT^;��uwc|ؠ��/y��,�m��+Ե,!�y�����K��FF�mlW�^B�����>�W߾�w.����8����"De'b��Xϕ(k�r����{�/s̅C1���E?��m`dh�S�H�I ��j�X2��F�G��w���P*0�F, ��nd��w�G���˴�M�\-1�L�|�0����!�t��L����,�;7rHh#�IZ�x$��z�Rr@�PٙK�Q<@f���"�ro.���m%&�\.�X.`|l�0���S2¡CG��,�fYW&
����p����,���Ln>�+y���3�`F����1~� .\��x0�Ç�ƃ�<	-���W�ZBJ�!�Y)���(.�#Y�+9�ɟ��F��nU
ʨT��K��F��U�0��@���'?�`|�����"n̼��w�?��/	�2�Wa+m|���7^��� ��Ӗ8 :�NA��
������WE�z��琥�gc#M��ԣhj�Ж��:�̥m��{���]Dƿ���?��y�{�R�	���(:�P���A���X��K��`D�t}2��&�
%��O�ۡ��5��"���a�G��G裨:̑_��&��B�J�#��z���r!�t��)p����0���Qk1�};*U�rR\�?jɭ�l�fU���bgxd�z��]&�F��H������NF^��Å
^�"���'����ކ?�� �9�[�A�m`�Ӽ�	.-� ~띿�FW_y�k��B��1�������<�2�#��w�Y�!�aU�gQɓ�(�c�ލ�{��F,dch0�n�����#{p�Z]Z �*GHPvX�g�n5�]H"-bdQ���h�3������ ��|��J�	�G#*Z��靖�)F�s��H�Y�Nt=e�ʪ�yl�������\��x�J�P�,��55����p����r�d��@"�#�}���(��%�m�1O�����m�����l�M	�j�(�� �!��#J#���8������U�e躉N�	d҇06~�/�z�BC�cau��X,���s�5
��F�Ƹ4�n����r��A�ZЂA�[�(\��ښ^�D�����`�D��"�A��y�d�dR�j �PXY�$ZP��yv�Z5%�šBI�ל�X.,��5V���i�i�.�kެ51{�
��Ed3a�N
1{��L����Ij����5k>X\�G#m�Ee�]9A� :<�bO�_�����gt鞓%��,v"
��fP+��[��3�����ݮj2�f��r���뫰iT�(XY]����S(���X���8��x<�maM�����t�d
��w���ԯ~�+E|멯B/ϢV���!���_��f��1~���k9h�j��L>bI����>�n��7.&�g(�`z�Xlj�)�y�M�GǨ*��� D.`��P�6?�z��#	zD�.L����9ïR��~�~�������1��߁��tIh�;m�/Rf)}n4uTJe�n�m�dV���^5�^�}�o���Hc�z��?��.���h6ېD?;�;��AF$��i�.�������ܖ�ٙ9�|y��|��cx�'`X
���k��"4�VTD,�Q�T��#��2J��Ӯcjj���&V7���� �����O�k�̬�w΢���j:�Tt��ُ�gt�K:N��2���S(����h)�~rW�Pdr���T�%7�t��կ �q;�)��E���9�Ff�k,P�Ty��{�l��,���H�p�gѧ�p�,2�n�tU��kkS�P<�!�d\S�>f
E�z��Q4t�B���{9	#	!H���ePH�W�����.i��@W��`d�	�&,��J9�N'MvVe$�QX�2��x���Dv �|� ��smh�鼏�?��\���[�����Ô]Hy���"�M
S��cj7!`ɡ՜���)϶L���P� �>�ţ����ۚ��~�{�++O%�������T�D�
$�(�'@��7���@�._��Q��V��"��_�j�T�O;��AX:i id����oW���E��H�a�^j���H��� h|ЗL�Nȱ\�bY��x�_��E�O�F��/كd��>f"�ܞ@�ji�H.[�|����
]�xb�,��5Xm�t�N��Za)�=t1������PБ+�� ��]�0������zѡ>,/��ā}�Mm�
k���n!�A��גx\�Ga�:�T��_E���F���Z����,KE�oD)��#b~i�t�D�jm�� �-M����}.L���),�O�/��`4�R�	A$G������uG���8a?VaW�b��V���H��S�ڕ��C�	��Fo��C9�cǭE��[�z�#hs��AI���k-	�`.�)�p�ô(T؏D\���0o��P4�U4�+���St���c�@2��]�k�8��U���9�Dj4�XD"jz ��[XhHM�D/V"��x<�q;�
�Ҽ���2I,��cddk�*v������)h����Jh!4��uK�~@��#R�m�!��0u�luGFY���{`μ�<��Y�a�:�[����5#pc����E�6�F�Q�(��Rc0D ��2�z���N� e ~�����M,<�;dP�t52�7;�	�s�����^Yz�Q�����F2�t6k�hC%֞�F`��tP!�F�#�1���>C����zT�*�A����۷oǍ��܈T-�0=��:9�}趽�0I��ty��O�w��~Mf��"k0��/C�AQ�4�lSEh�*>z<�����^ƫ�f1~�#8p��,LO�B$g����8��8��>��0����ON��j��P\C:�B�\D�/���u��?�;����x����`�6�����c�H&E�/���Q�(����?�.�8}�^���`4,��!��9��!�-��1���sm����R�"G�$A/���ihX�5���C'�%SAP���� w��@HU ��H���%���Я5p�� �?��;J��<���{�V�U]���4B# 1'�T�%{,[��[��f����zfl�ٱ�4�<(S�L�-Q� �H�s����ު�}�<���VUW߮�}�����{f21�NU�'��Ɖv+%]���bN�la�N;*��"�1@H����eu(��	���2��Gڌݞ����O����w8E<2BJ�W�\�F�ӥ�+��8�{?�r�Je�H�����N��>�VҾm�G�.�j'ȭ����?+֮��7�.C���Y�&Yh��[()J�z�)�Ӣ�+Nl�\�JY��p_t�����[����l�#��]߼�ݿ�+�³/~�1�'�p����H�,����,/穫�<��Sǹz�Ul����ERQuNFC>��_Q!u*1�وӪ6	�Dt�cz:��d��,^�����łBJ���4{؁0=�G�R�ɸP"�D#g���ı&�\I4�|�#�E"�z^��WW�)���mQ�u��؁[��X��[����<�ܷt�"E��1h�(9�����.V���h�񤭛�J���M��(�LN0哔$��/_�LfrL�w�Nӓ��UM�(��Z��� _��Gu�Q|��d 6���B�����K!+E��'��1)���I�1�"BqkK�]���?���8;U�l;�Cϒqt�j���˅�ue�"-)��1����z��b6�뱈ǂ�JА�3g�T�J�L������]S�&��:�M���}K��@���j̜�b�Ю�ƭ���&�>"DBBaYR+��ѣ���T\���#�(/Ù��u�Z^3�k۔n�����"�Qe~a�9ԛ��J��sDOק<1�QX�pbK�B��P����#��Yռժ�踎���5loW�Z���S�v[�p�r�I�2�dl$�oK�kbV��"�)�Q+la�D�)�&�:l�=L����[%���/=M���� O|?�+����}���eGE�`�B�!R�׫�&�@�Ja($��Ʉ�<����l�������I8���i1'-�Ȧ�I}-1�hRC�����ܖmr�#痃@I�]I�IE�m�L��,Pɘ���5~qzz��U�d�E,!�ϒ�	S�K2���D���SQ%؆_�W�YQ$R*�T���5Y�\WC�tkF3ì.���D07�rQ;��k���N2��	R���Cv�2��"wns�}�(K�C�>�Qc��s+�+��0�p���+�N�=ӳ�����j�Jz,Ö��3�^������%�ML��(�v��.ba���G���s������Ө���;wO�g�_t�!�ϱ�Y��/?�O�}��<��p��ޔID�@(�E����lV	���&[����uba��S�e����;I�7"$'�R/�u��L|�mq
x�%����U�41�~C>�e�G,��j�٦ 9��ay�y,z�Q�^�"�o���g 7J���eW�-��|r�TL?_ؐ~�+3d�m�.�`�rK�	��(����.�	?S걱��p:��@���3�bb0��*K,��{d�+�k� ����Qq�,�@i*���fQ�8CSޙ��}yS��?��-p�j$5&�Q�W�Uע�F���d���<r������x�W���~=�A:��O>��F��[+�-LO�=M"q�m�w���lHG��i�x����dBb�6h6�z{��[��^)8x�Ij�m^��q������
�z�H|P��f��b+Je�_�R"��۪3ݛ v��Pg�G6����an��}tZ!VW6�Q���'O(�Kƨ;��359K�i00��B�s�����	�H���4��u��>�k�q��tLX���6����Q�O\Y�e�d��x���S�����K���"#���h��ϭ���*�DP�EnSb�z�#�+[h�5��Y����*|
��E:*��NF�R���Dj ���v��f��2��_7yq�--�`K�-X!�7���b��q}�k��m否Vf(����������V�ą5�	�H���=S���5�z~m��R��ѫ69�of��ّ"�Ѯ��#����f����0�F#�>��ݮ&�!l[����m�;D6~�A��їhY�-q�K6��5��Rki�-?c)��-�۶���;e0�\��tz���X-�\�PR"�!�E�e�u�&y�";��Q*�:NOt�l�$dl�l`.�@����LX�vS�^�&�����'`c	�Q4��OG��j'Gb��ೡy��;��b�mL};t����#V^��� �6F���t�	���K���C~���Sf�pA����Jq&#.��S���d���#O��G����~gj}c������Q�'�xB;n��;s��ã:"��L�n����V�KR ��	�CCB����'�q%K(�n���v��&�T*-JlO�|������H�+����N�`nR��������^[�I佺��� ő���%52�.my|��e$=�f�@7є�Fq�po����n
k��G8|�#x3�`�|����kx������w��*�P@�n��"�?�0o������ԉgp�[���즚d���5mΜ���V�C���q��oy��hך�>�2'O|�����u�a���4�S���x�{�R��w�z�)\P��0�^
�^oT���?�R/�R̟#���V�be�`:�Z�N�?���r�Odp�V���h]��](m]'�+�w�I�z��@�ۦ��HB���L&�uB&�j��m��`J������jA�E(��uͶ=���*�Gu�Rjr�ȟ� ���[^AnI���U*����23�d�Y�gFuMz�,]�gc���G�7�SG��d�@��(;Pd͖���[�a�b��Xr���l}/bԳU��wC��D�(E���ĳ"�N�#��~&r?4��'��|�IQF��఺�{��}�ǟ�ߙ�����x���W�u��N����o��p�
��MZ���CLN��J�ӝ?���&��:uѾ�j��\
�K�Zbဦ�5��=#���+�L��zA4xU�[t	BTJu��mqn��X^;`)K܉�P_��v]|�A���_��"��������ؼ���@D�����@B�&;���nI����_����X�M��D@F��z�o���x,��f�R�x���$��ǹ}z��������L�d}���m��=;���S���).�Z��㶈ɨ�P��)9mڶ �C�q�4����T]W\�br�q�_�����Db�2�Ѱ R.\��Ĥ�\Tq��BS*tW�TC(S�V[�w)�M��aecS��2.�X<�g(&-:C��뫛��^�Ό���j:�{��u����h�m��<�����~���x�Kg���lȐVy�^���v-c��v0�H�'��(�z��g���oǴ�נd ��(�B��d*M�R��y�%���v��.�X~�z���II�ы*�V:U2�r�uQ�r���akw{��T�lQ�|a����)h=�l�r�Ffh�WU����pm���X\Gh�J��٥\�)�Z��V�I�+�c)�r+: �*��gILO��?~�v�$ݞ�gO�\^�Ѝ0��%�cE�ba��WQX�}� �c(3���[Ĵ!�q�-,����wbl���-
�"���虦�Lz���V��!E�ѕ$��.�R�I!,�_a�)�F�eccS%�g)V��m�ǉ.M���)*E�<�q�8n�j�����JHD"P,dqѿF���旘�>�Ӫa���4X��Z��`���eZ��4�"_)�J1S�]�2:4�:O�/J�(kVDR|�0����u-����%q94m��<��Gh!:v���i���_�~�8x��,,,������5����{����������ʹ�I�F۶�����(Ŋ�!ڭ�!�.����}��#׮��k��ߩWWص3��������8�|��p�z�����m_[��ç|�Tz��nl�A4�'6D�PΝ�k��E
�,3��|uS���]0��b;@4���3_R���b�j�Kļk;��49�=Mҏr0%'��t-khf0Fѭ�!�o�5ɸ۪�m�A���a��V�i�dZK�Y:��Wx�����"��g����+�:��E�:���A��5��tJ��l��Pz���+�E���1���	��(I[���pyq�G=%��.�"��u�Kd�8�u�,����o��b?��M���M��%qH��.3�hl�-JRt�c���>����t��ǆ�{7����7o|��
���P�&�O�͗k�o��:kUŲ���#۰}�]��T٦K����(m[7�r���F!_����w����a���`:LO��镩WB�~��0�^Z��`��� �Qn�n��]뉎K�CB,-- 蜮�`߾wp�}��}�y�̋�Y���6U8>33�/�p��i��N�*p ���_�ᨈ�e��׍�)����"�W1;le�hZ�NU3��+���w�u���L�󆕌/�Oc�Y'	s��y��,	���'@��gl�Qjf Ctv��3��>-�������U��/d�*	���:6>�`��ͭn���3ٌ�ha{M��J
�t\���8�R����X��0�1-�Dӗ��8M��\�Z[D������d�UZ����v`4��mTk[���e�Rׯ�h˫'h�-�L"��-�?�j�F��aq:[-�fE�D��ĥ�Sx�A�F�����_���DV�@`�y�C��.��ZϒJG�U.e����M� ^�NP�R_��ֈ����U�2�~��q:]���8�6��Y$�?�t�X<�I� �ZY�uAB;�Ⲽr�-�I0�'��S��Dv[�x�D�u
�u�Ô���e��>H�\c��+�Y����ꜚ��ն�>H�&M�^t��.�l��f+��4�d��#E����l�p@#G3z���e	�C:򒟛t���r��;�W�^ezzZ�߲ik�uOLL"�h�(�^?;5'M���XYF�ҥ�X:�ߏ=���J�@���kW�Rz��D)�7uľ������vǥ��x�.�J�V�K�'),p��    IDATl:xŌ`Y��ZhX>��F�6�V(ת�А.�d�v�DC!�il�t9��x�&����}��0D��������?��X�����{�����W���c��ۧ��t���;��� x��9&�}�y^�Bv�H§��\��a�x5�W��A��y�g?D�ӣP,��x�����gٽc����U_������N���3:�7�Fƶ�ǞJ�N��Qځ��e|�I&hT6�o�cx@ʳ
�R�rQW)2#�X��)�&������h�Onc���O�nc�Pg_�Qs��{�L��z�s٬H���Q%��������ۏ���9��H�QY�ϟ����=�H�Xi�r#yD�+E�6@jh7���y�"$R��9���&~��`�C1�,�޾���Q�6����Rl�tHc�k�`��^��ȓ$�D�j7R��K�ZI鮋(J�"�ꏊ��j�oޘ�����s�Q"��JI��v��^z��O���?z�h��
�7��:��7����-�M]�kVX�b�\�C�����$*�i�2�ah^�,6��N���&�25����I����|��M���5���x���"��2�;$�70&m0�M�ӫ�M�7��$�]�H֯�`��ٹ�~N_�׈�`�da~Ík�i��>�P|����P����Rd���XF�z��pjAsTkm2����m���j�L$��q�_\*sy�ΝoyG��.�++x#	���#��&�Y�)_�i�x������-��c�4���?��%ҭ�1;>��H�6�z/���8�
�Ӹ1:鋟�#�Z��e���n�0�D�1;ll.��p�˗/�
E�&�%��Tu����EWn��*<�ݒB��c�F���?����T$�.��x	�6�W!���&��yQ;;1A�x<$bIv��҄�C���t�m�dJ�^�,�Z�F~�+�N���gמ��=z7�F��Gȩ�տ<2v�7!@aq^ouac���;�<����Z����{8���N������V��vK��u�[Cc�1�檘�K�O���?�Z]V@v�/�C�щA�����2��,^�g(>�W�Mb^�\pkR!���7�x��O��zZsb�U)U��f�Z�(s�m<���k��&�IW;W�,^>��FB�I���|���F_ D@�%CC���S7���O��+'�`z�v�$qg�y�'O�i�ٱc��3���?�=�z7/?��ܜ��>��];8y�U���8y�$��\�ȑ��ܹS&�B���O?��
��+�_��'^9ɱcǴc(����|�#�;w�����!��ƴ:�q׽�����^�ܩ�yz���T���Y�-W��Ο=�T�{�<Q�Ѥb}��_&�r�Ȏ��0}!��/q��^�{�fM��L����Ҫ:��f�j1�i=ሏV����:#�)fvl��?��؎�s��SOr��	�0��6�������w����l�c|�v�K�5x�;�M(�K�0�sY�NW���b� [�,u������P�Ui�m�v�������괖.�3O��L4 ��6��5<�$���Q*��������"�dse�������������xXdkx�t��wǃ\<�cd�V�����>N98�����H&��"���X�Z~�V�*��"���,r���L��p
K,.���FI	��\�V�`�1l��Ǒ.�"��}=��Y-��b�p	EN��\��"W�5G� ���} 囹­�z>6�l{�hb�X*��|x�N�N���)\S��~��-�v�p0��)�x����`3_dy}C��pG���F#���?SRS$mŰu�|3®_J�*�I��P�5ȕ�����%u�o�M,AW��BPM����H�6S�d�O��͟~�S�Fy�z��������+_�J�|�!��Ԏ�����R����!W�+���b�����"6�7@�TR7�2	��z����G�4�M�(۶�9u,�������p"܀H�LR�qu[f�����!#	9�E���^2b�8sio"D��K�n3əg�>cl�`y�9V��R�m���$����h�O$�\(3�w7��5�ʈSt!�F��&��-^��If�w�� �4�M�))���Z�@����מ�G�<�P���G�V�lt���qLa�	*���LZq��̤+#DS�?�&���-%�ډQ2�+A��;60,?_��գTZ���s\�rFSQ�[G�'2$ScD�C8�O�  �uY�JZ��Y�چ��\�\�#���R���S�*��z�H����ܫr��Jh����8����Ro��C]�-�?v70� ���]���+gY�\��c��[U�e��$���.XK���a���%D	9u4Z�^)+�N�#Ã�on��n��^ƶMSot(��W�m��O�ҁ���욚�,]�.�r����v��s'��JO�*��e,n�T�&����h��E4-�c� ��"�jk�5D3T�_���9^=�M���x:e"~�͕,��'D�,ƉA*�M,w��<B��ei��r��r�D�m�HMq�������ɉi-�~���������� �>��j��(�����U�(E�]�?�3Ͽ��|�����/�?�s�OO�v�6D�(�g_x�\���|�A�����{��?��)^=uBu$3�K_zLM-����y��G���߷�����Hw����o8����;�����El`���?�3��ܟ����|��k����p����O262������>���8�H�W_~�f~E�w���$�]Y$IP�����i7*�z�N�v7g殩l �|���O�L�D�YCl ����G�؇�K$f��s������@���k���O��[��_}��V���(咤,Ey��o!�TN� �JkK�֗9���_��#>���)��#�*]��!�f�R�:�_[��3O�Ņ�$�DB2��°"��~�p|�����YvL�'�`t|�/�>W&S!eΊ�f��+d�@�)16������,�Z�����%�5r�BS��1����K���Q�^s�͹`���{����h��v�(�W��TA�<N=�����^�z<t-?-WRU��,�~_� R�v��#k�O�/�`q�^\G��Bq�Q�E�b�&W1س[ذyl�%�w�X�J���q��bX��tǱ�8]l�pj�4�=.__�"����f�έ�7{]�:��Bдxj��Pr��δ���.c�n�*lk��E����E��!������bϥ��JJ��{�����E��-��x��*
�����;���ի7��:>S6��&}�A��cP�fL;D��ֱa�\ӛ��R�H��8��$��!�jm�[&�LQ)ɍ�%�u���.�%#��Kǒ�'E/���)d��i��x\CsL9�h�0|�x#�hY|�8r�][%-����D@����w������U�OM�ml;'O� ���EO$ū�q)TrD�!�n��u�P�c/�D8���J���{/C�����e}}���E�!�&$�í��L'�۳���yV���k��<�+�z%���c3�Pk�s;}}1���u�N�e)��p�D�&n;��
ѿ'	""u1����x4�C��Z�W�^���)��by#����,�@0�?M��Im%�>5�|��xPW��pX���O����R���܎��e"jR�])��ф�mE��tmҏ��ו���*q�k������Eq���۳��bx�Z펪u� ހE�^�� `�{*�3Y�E����((�YJ^jG�ߖ�@�WV7�x��2��K!݈���:f�\^�xC�qX^\b0�b����e.^���7��o~�5�&�ՐRn�T�(2�J�xع#C:c��r��x�_F�1'M޲b�矧^�Fq�$�� ��A��`%�ٮƓ�_z�����v�|�8��\���9�_�np�Z�@8��_�"��O�}�.v���W��8������!���w��[҂!����������^��=�mw�G��08���o>���"��MvLoW����H�o<�-�=�G��;y��+��_�E���/�������СC�������.]�/��/YZ\ֱ�c_�2�33Tr9~�w~��~����q�}����oY^/�����׾��t�==�����kE��+<���l?�g���8��q7����>�e�%�v��g_P#���|��>E�����~�����mx�30���箑LD�-]`u�5��il���o2=���n>����48{�9r�yJ�<�k�$�-$�~�]������?���&�p���!�d����;�_;�W��Fv��W�����=G�PY��Q;�ϖȌ�"4���\����48���h7]�j�c�D�������"<����>��O�s�Qb���ꪷG�q~l��/����l0�}������课N�g�]�b��µ3��I5�"��$�0�b�׹~�	�s���ﾏ�����ϒ;�$�DR��v���Nv�4r垶�xC1�z?���S�IUb#mS'H��	`^�Ҭ�_�� �Daʺ'HY�*�����X+4uѩWq�^����I����sV����x�j�HW0Y�(u=^W׵�i�k:���Ӥ"?�e�t�++����I��(ES�S[���W�;��6Ȟ�;��,�J�]WiM��j�0<0D�����[��qߟ�Q�Qܽ�+��ǿ��fu�a�סZ���5��\_�E���p�q�e�V�QB� H���&Mi	����m�����hQw7�%���3� �vCƟ���CU4�!����2�!�ڮ�F[r��::�bEvu��Ðq�gt�!Zf��N��w=����h�b<�	�������?J4�cthP3p��G9u�%*���jJDMz�)(v���Y\'�O�?�/����(U�,�ɤ��EST�y�J<Xz0�V��������m=��Y�<G��J&�껖�\�Y���1_? �
��R)�\�����O9���	��4�՘'q�J�O4l�@:�Β���#d�]�CA-���(#-q07���W��`�4ܺ�p��'��ҭ��%ڿ��3��J�&K�>�� by�)�Ҿ>F#Xa:8���aG4���t"U� �#S�ʚv"F����p���+SSW�����kv5Lݚh�T���%�ZP�%BO��ı"Xy�"w\}-�?$k��w�j<x�x�g��x��!�9�]�glt��aVsw-O�x"%�b5��VR?�� ����;ƣ,��
�@���� ��2�HG�I����#�{	�t�\�t���+x��z�W7Y�W(�ی�o#�H�cPڪc���:Q.\Z��8wu��2-�d��a~���d|b�f���>����W�N�������y�xD��Q�S�������������wPQ3���?�o>���7�z���
�~�ԫ����Խ{�Mw�~��J��y�����G?G(�C��v�s��i��o�V�n���ԧ>����f���~�����!~�c�?��,�Wt�����/��ػ�G��2#cd�V���g|v�w��=�v�[Uk��Y��'>F:�h7�w���}�Y\�r��1�����ӂw��g��p�(��5�����8T����w���s`�Anݿ���~L��@ f�Z����&��S΃�����|���ċ�?��3�=�K��-�)T~��=p�
K��y9�����E��ϕ���l���M_��^�K;ܫ+�<��o��3����&�z����oH��_�.��	$���)�s^_ @��N*S��H�����k�ص� �Wm�>q���|#�)��'����0�#�
�vZt$�^!`�	���������P\�H��w	Z%�d�zG�q�raM��Y�ߕp�.�X��{��f�,{�8�e�����'lRq΋6�����v���E'�-����̯e)�J�8�Q�ktiɽ�R�~(ԣ�qz�<|�Du뫫�X��[9����e��HЏ�6F�E���T}��d��]��jBݑ��K��Rkw��(H���a,��S+2�]˜Ӧ�v�(�������y����}�z+�7����4�)<��_i�/���2j�ߨ��N�t�Hܙ7Ln�A�ܤ��312�����$�U�_bnЁ`G\��� #��֛:�H���9��*�b��HHڂ�b|8�z4�L����Vy���&�Feu���5���C��O2��ʎ=��p����%p;9^=�=r�W�f�002H<%"ܵ�"��K��^��I*��[��8�����������޽TD ���F�W�H���m�����E�F��x�<��:��#lT*����+�V6�61�ן��;�arlP5��p\ǔA�H籟�$4醉.O�=u�г�t��%BpɈ��(I�f����%Q�����A8-��I�ev����	�ڃ������H�.�G�v7c@��%5�lH=�)���b��c+4	�+)8�7'h{��h/��n�����g{���%���v��nS���T1���\ދ,����
ӽ��J��\E�K�&"Qu-�.���Gxzr��vfpX;�x�P<�,D��$_,jg빟<ϱc�u�g׬j�^=}L��햡.�[nݫ��b����[�%-���� ҫ�~�y�w��;$�#��k�e�v[>�)��{8�f�nQ_z����8�"�D�N0D��%_hi�K�N�&w�k�-���]ɳ�-q~�[���<��.��[�s�dǘ�����k��kg������ /<��hCA~��&32J�Z�_��O]�C���ȭ��F��O~��b��z�-�;x��B�,��K?���U�� {v�fj|B�i��Kǎ���l��{�t:�)
�]�U���A"�(�@Bƫ�)CR�SS3�=��)��=s���.f"=Νw�O�Z���>��J���w3wy��ɝ�S-�_�������{H�X����AOWe�~��^����I��<��A5Ҝ��H����Yݬ���;~�o~�{|㫟g �$�
$�ή����z��Ѥ��d��9fSD,)"zģ)jWs�-�E8�鶨J�o�`rC�I�^����H�F���'��bht����O�h��_}^������ &�V`�P�o�]Z��N?V�X_x���k�L��3{�g_Z��/]����Ij�-�w��ٹUf�O�3�pn$E�C�_�Be�$�|�r�ѽ��}&{��K��箪�'�I�A��,�������d�ꌮ���}��U^������^�a�:"#c�jR53X2���Q���rz~��>�6��93N��SCKȎ�m��4�*x3���ē^*�-��z6����%��&�@�l��=��h^%ť]/���,�V�����9S��B�
fF$�NǠճ�^��4y����m�l��uxj�&O�B�M85H��O���om�ԟ<�?�V�(t޸�W�uu
W羜�x鉿o��:�sĢi��+]�N��:��o@��/�	�Fs��U���ޮ�զ�4U�.F�ˆnң^W8m��ҵ�ΘےPya���� ��OQ2)ȗ��.Qp��J����(���P�G8x���1{7���o�p��9{�*���bO��ps��+������62� N#=l��V�	�8��ԶƆg����7^ +���,�f�|��w��6�=��ghdo ����q��}������g9��v�=���Ɂ8{��p�-{U+��1�\,Ke�\Kc6����T��������?���~�%�����%�q)�ndo��^�1�?^S
5�ovof�����!������H�O᷽�>�Uޯǃ��_WN��|K�ǚ�F�n��'~9���[t��)�Q��[��Ot��ϐ8��L$:y�8���5E�#��äݐ�B@��e��*�L�K�}����c�m��������_Ӏ��55<����p����\�A[*��ַ��{����e����H0eǮ��(�G��R.�ًgعs~��m�q�#�Ya�Nw�c�Se Ӎh��9��=����	/<K�W��(��"4���z�`$b�2㚨R�rh��x)��;sB�^/<�#hd�onR��aj,���ܞ���
q�k�Y�j���n��K�Ж}հ)�2C�4+5&��Jy��!�FT���\e��$�f�j�F�ob�}lUĸ�~�P�    IDAT�=�acE�4��緈�Gi��,_/180���:����];YZ^Px�Pd{2�.ْѢ�l�����g03�H�խMv�TlQyk��pRSL|"10]*��2���۰0�J��il�%S�T(��j���������<���;9y�)��E޴=��Y �ORwLέl�P��R��S���#��s����?��] L$2��mG�,�1��v���a,�]��h��%�����?��s��q"��ΰ�Z�w��F�(S�H�@�Vm���I���O�v�<�����z��T�\��'O���}�k�V7}�P�]ˑ�8N*�bx@��t����C�n9�]����$F �Wt��2���k��$�~��������g���!���d��3��?"(��:�'� �L�ڪ���TKu�}c!���ރ���F�.�>ڔn���c�v$����W�塐�ѭЬW5+=[nS��Ć&�L��$�
a��¿+9�_NQ*m`�y��2w�DԏS׋A�+�O&�X��:��n�~8�Nj
��0�g!�����,S�n��C���gyo����Ø��@8�#�B����v���k��uM�e�R&���u�C�������7���U���]��U^�����~�Y�{��s(6�c&"�j����m��W"�$�@慢]�΋l���aө�̤(��ZT�b�6[���}�t�����n��p2��}:
lvJl�slek��VK:f$F�k0��]]"X�I�tχٹ�>��/�j����2�����`�D�B��ɶ�x���_��_�k��W��]%�����Q��g��,��A��͓�MU
�t2��0Y[Y�k�t�F�d*��Ɨ/�iW�fRÝw�����~FG�5�X
,y��8U�ҏ>
�D6I2���}�P�5VI�7Etm�>S�m\���tؤ��;u7��v��xɿ�y^r*�\n��X���'���x:y\��j�;��Z:�����W���]Wߛt5��SH���E���+���iQ�V��Ct�U&�,�7�n���������}�b~�W�:��w�� "t{�Z�s�#��Q�o��+��N�����y��cj�����T>��(���78z�vu#^����O����8�^d�����ߵK��յ9�v��oϰ}R4S"̭��8=�ae�J��ah�#�����=I�]dp H��R*wٵ�v
�*yӡ�(¨U�F�M��P�6iu{̯g��w�E��/|z?m����d��|b|�N5�Z?;4�4������K���#�F��s��\�bE��G�����#�VVXX�Rs����ٍ���h�X�78u颀��4��"�߻fYϖy��+��.�J������A�Z�B(Ҏ�D�M������c\.��9E�Ц�Z8��r���+����p<̘���]�j>}�8��(4�,\��f��Z�x(�@&��s��3=���h�U�|ia�+ׯ�mj_x��]��h׸p����^�������r���yN/ey�/�
ci��/�)s��c����vQPL�=jV9����?6Bik���M$'/љ������/�����p����s0{y�\=�Rv��34���I���Z-����O3w�2w����Mau-�._#�ؔ*9��֪�sk��3	��=��%�U7$�m������F��*�h`H�u�&����Z��?��t��q>�я�r�E:�?`(^�ի`��c*[U�V�\��_8�6[��H_L��5�tb���C1~U|������5�	ЩaQT}�����c�3t<�=��-:�f���E5��^�ݪc%:�&���ou��D �f��F�01[��6Ctt]�hV)DC�zr���je�4:�:�ez gnᩊ���f�5ק������A4���$Y�
��C�)
�Xr�z;�M��+G��ÿx^�F��z���.
��}��v��}X��\V~���r+�F
u5o�i�i��dҺ�J,P��bߎ�����8�C���M&�.y�d����{m�n����#�z��^^�g=��בS��z�U�@4 l�$l��B���r��v��~��~�+YW7��[�%1L^���$FR�	{�G?�Qd��癿|�\�5�)S[��b���0����b��>�
ke����f�+7�A �^���8��G��;k��؋,,\�{����8?��.���_�x�h!�S�=�
�ear[-�҆S��`M�F�'�ą�e���e2+�K��Sf׍d)�n��@����?�fR����E�jvL�.X������S�����b/���??������4'�¬��_X��l���YR��ߛ�~������o|ݛ��\?yn�{�_t���|��zX��^�B;&�#�~t�l<�W
F�Sa��h$\(�M@���X��y5|�� �+h���Sz�پ}FcG�dcn(�e���f�\.ˮ�IFA
g�-��I�ƽ�|M2鐤'+�)_��M�bt�=Gfh�����'�뱹1'��"M�"-ʝ5Ɏum�A^i�lt�Y/5���g��b#>�-�kBE�i���\�dtp�z��ёk������S1��Pd��V��E6�UB�������	Z=�
����%N�=Ǯ]�ٳc�Va�D"��F�S�͓c��E�=���ߣ]�|��Kg^��iW��q�h:��z�0�Z��Ɂ�mڝye�*��r�����c����*P���>3���u�F��o9��@�g���f�D�����s|t�=<�I��X�"���st��du��6����=��	@�f���b="��Q�1|��Z��&�9.?<u��zϿf|�;�re��}�O�X>ˮ�S���F��圚��5(om��A�B���I�ebX^��Q����z�Ȯ�{HX]<�ĐI0d��+f-W"���[��QR�4���p�̫��yP���)ӫq�2�m���tہ�X[��u�Q��m�x�6�y�<�L���6��$�V�@tZY��Kg�\�­{���r���'(l�S+����m|�c�dy����"�Pi��-L��v�d��,^[`zh���mm��q��ܢV�Z�M�Tw��Õ��_�<���_��F��L"��gui���aֶ�j�K$�u�H��4�8���w�v,�8FϤY+��*C�:m"�(�R�+R��(k��Lbt��L䎂��2�������t��]a0z�((7[M+"A�����]��!�Fϥf�(4ۊ��Z�Nf��O����ꍢ���Do<�u���?�x�r�>�+���B�yjҖ��u��Փ�Y;�#���l?"�kR��m�V�K�?H	[/�|ې���=�m�Ѫ�-#�v����Go=��3�Qm����;����i4[!E��A2�#�n��a&�;��ed�r�*�_?�+g�1� ���n�D���Cw��ߢqs�n?Jjh��WO�qt�kj ��
�-d�4�Q���ur6-���_�i]��l���
�g�O�y��6�Ξ%�]c}sM1��?�'�ª�K��-A�wnSP�2Judl�G-Ȣb���E%�G�f�z�Z���E�$�7G�R�I'E����e�!7)���ﺺ1��S
-u�z���`���?ҾQ����z(0-��}���k)�_r;���/:�9�A}����5��'�F�E�ߥ0TPy���By�5�z�Y�, o��s�c)�-�U^_~�MGZ)3��Z�bU\��i	S����'���8���p$���p(F�Z�$�~qx�'�x�����������j\����^_`vvV���F�F�Ѥ�i�.��ؘ#df�m���&|ʭLDc1�]�l=Ȟ�"�m/��/��+�bz���(Ӕh��vD�ѡ�7h����D����� 2��'��%�5�p���2��T�
3T�auM�n�X�C0��4���?K��	��\��`�P׃�覆��S|��3W6٪u�x�;vN23=��������-^>}�Pr�����γs��Lo��K�O���E&6M�T&�P�4�%�p<���]��fiq�ӫ����y�������K0�Z�3�I�ٌǃ��\�v�gϳm�.J�&M)0�gS!�nM	O�ɛ��crp���RCc����fӖ��0A���҇2A�^���;���HW-H�����Pr�� S��l������,\>�-{'��K�}�t|�s�i�xS��V�	�-��JB��b�Ex(L>[�n@*5�r�D,%�01�[[����J���M&w����}�������{�Iz�g���9Ǯ��=ӓ�f�ь�(�"B�066l|���>������`c�9�$�@	��fF�CO�\]9�t���4�.>�������ꭷު������N���~���v��ͭ�ow8���,6K�Tl	MEb���i,�6��Mt�ίq��iܾ0����_��C�Ґ��f�o}���u:֗�`25X^��ց���w��WOR��	K�ZGj<��"Dn���['�N�R��bbT���㊐/k��Z�6�6�Z�&��NU��5r����\G�v�
��r�_�.v��i�>;�n�r=�R��յ,D��!��y4�"�V�Ѫ��g�5W©Ef"z�rMX�^��|5ju9%Ww;�(���V������S�y�լ1+]��Y�Nit-�-Y�ĥ��S��Uc�X>���h����G>�u�����up�Z��k����.^��4*���tuU#�:��8=UӇ�1a0X�x9���$Yp��php��j�J���,,-(3�|H;����6��E��j�I�ũ)��V���Rڎ��2ѡ~��h�-���Q��#��'��&������>�Y�����n<v�b���<�w;��K<6Ǯ#�c�.ՙ)�.���-#�xB::/������������<�_ؠ�(P��$����/��絫q�^�pI�&|�ӟ�{��h���nְ�j$*-%��O�,Cr;9�6���t�J�E\��"�h���vFfŌ��A�1���P�rY*��2�"$����^�E�Y`%Y`2�Rܚ�\�W�'��'b��Q���>f2�� e&��PU=��:n0����"]ѽ� (�S��T�vV��LJk�F��(ݷ���r�i��lʾ�J+��56~�$��= ,��m5���h�l�^M`�&��F|���qOG���Hʽq�����@��@N1�w��_����r�z�a6o�Ɨ��>�����ٴi6��'_eמ��u*�.S��K/r�� �}M���U�^�aS@�.,������3h�����,?�QW���(ES�V�g@�i�]�:��j�jK��CL/g�����1�^hap���L*�HB'�/'�Y���)g�t���d:];�kMfWJ�n�n|v-;�8�:%�/ջĲ.^]`�֭��з2�*e�U�//RhjH%�Zn<��n��7�be]�[4J��N������^,N��K�J[CU�^��.�;�"���X�%z��6���L$�&�h��*��5Qi4Y^_a`0�Z�*�.>��(]�),:-;G6ch��ܕ�������\��m�Lg���]V�R���ӬaK$����fh)#�J����S3��枠Q����R�2����t���Xʦ�Y[g.���tb1X�W*�ő��`�k	���*q倍��j�� WN���vsh�0�|��v����Aru-f����)�}���(�n�H�.��)wh����D��H2w�<~���v`wKV��a���ɖ�<���hjE��՚wp�/���v��?B&�́-;X_^$�����ٖ���_2'9s���8)�V9�o)M�d�vu-�o�۩kDJd6�*d�{�:v�E�zq�<X,�}.Q��h��4K�3.:�*�n���4�ق4ܸ�M�+-4��m�5e�Tr%CQʙ2����ɱ�K��k*�����ؕԃ�*^h	3(�����YM�&1��`U'��JGM�v3V�E���h5�UO{o���M�Jz#�.Z��:%}��V����v�"�G>������~�׏�k�g�|�;���Q�]�F,�S'g>��P,������^Y�Ę�Vu�+H��K���>5Z��2�
�����:J+ҬV����L&��.ހ���i���B�z�����B�J�@0����(�\��%����j���KC涻?��=©�gx�87�@���q:�c�Y-�o��>3�f�}��@d����9y�)��%4���Y�[X�k��.h��l�$�:��a�P�3Mܸ�!NB�iR��_~E���?�5�=��fS�VL6����E2�����)`o�	�Ql`Wƶ=P$�TJ���H��k�^V��n�2���������wa�dl� ӯL*=p��
[)ao���*ӈFd����i ����>:�Z�}U�Y�R.R�h��"`6�%d���;����kf���q�;�Mi��T�6�:*Lδ[-��-��5�`,�^�
\��dd�P��<��B)�#�H�f���xH�q�\.���M�7i���"��eu���?���_��{/_��������jQ��AU��+3��]|�26d\��a���4�z�̤�+� � ���c�n���=�m��"~�V�4�j�[�P�
1N��8�n�&q�k�h���~����z�|Ä��em}���A�ci�� �_�ϙ�Os��ǹ�`��F�Х�1��RE�t��F�g#�>���bh��|2RNUh�`p��R&N$h#�2G����q�}c���.�cl0��aau�2��Ī<C�ڐ2:��M��]������GKm���.r�j��TJx���4>G�j[���wqʉV��AƱ�:��R�(��6�uT�K���7x��o�is�r6�hd�����0��d�&����u�$�)��6a/�\�_<�c���h������hȊ]WQk��R�';�.���o�Z:�ْ��x���#:U��#�����
�
3Ә�ұZ����d]X��d������1��z��G�pЂ�e˞�:Fк��9���&"�~^��Y�r���U��*�bIu��6Z���A���B����au������l,Ėɦ�g��VS�3�/]�3<��+��h'�`i݌�n���2�����K-]$=�*��'0k�1�5*ި�p�(�I��Ũ5)V���L��e=����0�N��#��"�Q�t&Z����T�n�!�8鵖�jMV5Y�Y�*-@:�\�ˉZ�S�c���6��F1��SG׭c���J�c��?ȸ��͖uU�u�}-GR&k�N׋�9�����R�@9�ԫ�;�[�����b�Ѯ��4hv%�_�ZZ$z'%y����9Cʖfd��?�����:�y���#�k���}�R�T��XJc1
 1mX��R@�T���tq��Ŵ�utZ3�t�N����/T��=��X��>?�@�x
�ΠƢ�R�L9�j.��?HZ��&#��V����ru���W����zNse#um����0�&�c��e>��/���=�[�Y�Q����H��C� Y�����?�Oy-�g��c�-E|!��
((U�t�NV�Tj."{X^�357�u(y_��c8�����y�������7�<z[/#��P�p�?��cjd*`�Ѩ�3Yx�^�b��m�^~_�����F���1���=B��
n.ĵ�+= �S�k��m�Z/0Z�wM��V��ER�{�Au{��Uzc�ޘ�ӻ���W�X��NF״�z���h�$x[�I/+0ً�O�Fy�:C�6�frFZ�4����F�KmTӪ�z�_�O@7�������-��V��W+�_�'7��!W�*��ca�-�3i����ϫF��;w_]Ul��?�9.\�C7����|��*���7�?����!���"vM��p�5�H��A2�t����Eo���3����;�\|���W�z�^`&���i���R���0�tXXϖ�[�L\w'��a*�&���M��a5�L��N4���Yo�
?aF�u�g)��"����;�����n`�����⹗٨��q��ή׺���!���b��M�34U��Z.���$]m��׹q�-�W	�#hz�+��G�p��	���l�;7��0ŊM����e���E��u�TV�L*�u%cfy�$$_�hDԯ�極u�n7�v�D.���y� QF]�+|�_>N�g���pˑ9|�=*�R:����V��%    IDAT�дX�/�0
�l�U�$?��7�c�
�ܲ�^=����_���mߎ�7���瞻�C�(c�k�xa�rGG	=f_H�9�^�/_:Mb��^ �R�-z㊘��5�G��6��9����aq��A���7������O�S��\Ř�1w�$��5Z4X-dИڸ�:v����}���m��#[M�(�Y�\9�2����;5�N�������4���`��0؝l��f���P��@n���ǰh�t���*퓢ÓL@��up�܊�-�t�ֻm
M=���Q���,,�	xt:���YHa�kTۥNk��5����J���8�N�>���M]��ꔈ%9�֣i��w�XuYt]�O���I���H	|͠���=	�A��(]�	��`V�fa�%�L�lY���5��p�2V+b�ͬQt��q�CU�Y�H�۠e�Q�����v7�CG?����|����o��xM�pm�'�Ǿ��ja��ҤV/(P(�R�Ey�H���a�r�V��Nv��JY�|R]�����ܠ\�хHfV6�p� �D���K�Zarq�X!��e��i��9I����ؽu{�Ӡg)����,F�V]�_�x�x�Ç���O<�c�=��1��b����d�������>���Y�o����pjM<���ɖ��꫘-z5ڌ��C�E��O�����乫dkU&�oS"eѽYu�f��>��c�߿�-n�����2��(�R.� d��FM���������i�Է�J��|	V�W�/-@�7�U��\�����x"�!�F�����3�F6'�*[PN�eF�qs���^�n�%�ZC��J��<�$�PrEG���	dt- R�Vyw^�z]H��,���M+��.��\��J;��5��b��(W�͍�/٦,��N
��_�S����Fَ����jS�b�TQr&��l9��z� {�kZ*�B���ڕ��Ivlݦ��ZO�|UEм��U��Ͽ�ƅ%�/���x������P��7����2��E\�{��{���=�Kv�1�MtfrMێ��#@u�<O��8te�"v��&��Y�L �t��{�N�Ц�dd���;��&6��|�QV�9�!F�*T�54x�n�����HN�YGj�,�>�]�F'�;ތd��(.]���'�3��1qc�5�[��$v��c˾�i���ְ03KbuQi�����?I�^�f�1�7ƞm70݆�f�S[d���{�Y�����q��C�J���~�����Y��q��aR	{�	u�*�\1���b0(��¼�ֻp:͜8��ϝ�l�bq�y�o�!Ao���e~��/�Iϫ����_�Gk�S\�Q�4�w��m.M]����������nbj�vS�ny��[��>P�&K����WV�L콙��<۷�`߶	�u��1��f����X|~�Z#w��f�(2{���fb�38�v��&6�t��|<���7�t�g�}���Pt�f�I 4ʅ�9̮1���_��,Q�шTEF��L^8M_4@�:�F�N���`"������|���2LSc�ҩ�<{�A����23��H���A�S���x�~��~
R��ҷ�&4M���)r��)���V1�4�5�܊Yb\4�z�I��7:��^��Z�K���l�ԉ|9N�]D�iP/e�h���\)V�k�M�bא�%���T�-�l�7{H�8�CXlaJ�&m�Jn	�-O�GCY�u��J��6��C���}r��Z�D��c/�U2%�G��2�1Z-�gV)�
��.<NwO�(�z3%a0��K��$	:�&�BU `�Z������4�o}���~�#�@a,�������J��&ɡj�T�����>���$�ʫ.M�3��R(�r��?�tk���֗	��$b�&�Z��[Y\"���/�I��L.��2멙��,�خv:�szU�rl��x�B�J��0�&�iiD��
�F����!���{���\�Nb6�T(�Ӫ%�~�_>��Q#��z����ٓ�
��꥿8�X=�/B��dv������~*��;��2�I�ƨ�$�����s��/<���r��+�۵�n�����`!�g��m
����h���� ��O1�;�z�7�7h�Jq��]��

P��~�'��Tg���2)��26���`V�]���!���6'�lJ훌u7�vUE��;��Q�7a8�ofr�+�Da3�	��'�J�'�MF��l^ݿ�.�M@��D���\�3�%�Xr�8m0�
K��5�d#�F�C����-�V�M��>1�H��P0�~|A�mN{/d[�m[\��7P(�9Op��	�o9#�K���˗���њ-L]��������X���?��,-��&�ƪo�\���B�&��-��	Ơê�b0�)	ضE�~�=`q�˟~���a���׌=�a�~J��M�W��z'u���.����}�_>s����d�7>�:�gϼ@t ������o����Fxh�<���s��0�m��+v~�N�O���S̉�#L���-��ի
3t�%9��+x#Q�{�C�JR���L���<�.�Bx$����l���M�t�9xzC�����+�ii�}��L��t��=��V�v1ˍ��h�u��zY�ty}Z�6R�C�gΜ!��p�ͷ0d~���ZC�W���y�o�DG��p�g���Z�������]}t�y.]8Il}	�?�����/'�36:L�T$��L���a�eԏ߮�e��+u秗��a%��w�ϥ�W��̄�>�ٳg�:�{�t1�����G�w[�;���)��5�4Ү�hw�T��<k���ea��m�rL��j��M���D&�ej�4���l�#}�rqe�t
t�j���Z��.��=��s �sO<��8MF\v�z力%r�4[��)�N�\èӑ�'�^I�����{��j�_��<��g0��0�eAM�Ĺ���T���%�:wU�����*T�B�����Ch�j����4�X�lT�[/c��1$
m]�K���[R��*Qj#m%��c7X1��x-5��$�nY�o=�M���&Yz�%aAj :�Ɍ�cI����#E�^K�'�e��k��PN����jҦ+�&�5,�=��혌��i���k���&mP�g(�{�v������k
-X��}��
ϼ���U�Wo����r��T�E��%�{�$IE���v�>�fNW�|���ܢ/:��7�U�d��	L�:n��t|	i.s��,v������e��0''/�V.yДRڵ��A��$�I1���4#�|��EQ�A���#�S�vɮ�2�u/�o{;��J��J��F)}�_<����ߏի�\,�5z�٭h�%RI�&vP��0XL�fX���^��,�8������rB�;�
��%������|�'�p���X]�!�K13=�@������l�',U{=����\�N�ZQ@K`�-@K�2Ѧ�m���0]���0t��w�AT�k�I�L����]*�����V1���}�{T@�H�#�G;1f��J��t* ���///*`& P�e��#�θ��l��~�XV��d����n0�9������$��Z-�s�|ҋ��+�&�M�ܲo�0��=糀	��v9ܿr\�~F�}J(ב5����W�&֗�x�g�F�>|HYY��6O��J�2j�,�a$!������TYh�c#8�ZbK�.�捷LtWp�k8L:U�e��$m�!q�r7F���~�2��0{�5��C�q�u�u�5��p��o:ȚG��r�Z�����'#=2��F�@�&5��^fߎ����ꙧ�t*lں��/>O%�H��'��n��&��_"��bt�^�r��bBK��"�\�lipe�s������X9t�N�m'���8x�:r�]c�=��[���ɨz���z�ud�晙:͙K����bہ�LN-��S?��Y� 'M�~����������~����h3r��y,����e۞=���M�P��_�'$��1j5#c����w�67�W��6�;Ԛu����̝y�V3��DT5��ƫ\�<��-8�2�4HC��F%������ou�J[EGC0�O�\#�.��{lչ-�+�l�2H�U�PMS,�yۛ?�p��'�U��"��b6�A'�vU�נmR���9�|^�W�B��R���t����X�7�����n�������=>^�œ�9���
�<L�ۤZ)�-�pY�k�������G�[X�_���#�i)�Jq��Ef�8z��.�e� �'&XY�cj�"g.^��v�����j�?���q��$�F��M�X�$l`���WE$5�a�$�(�/ښ��D�d�mp��;iH�A�����b0�OK-_�N��J�4􆒪�+64&lf/Z����K�R�&���AW�Z&̀O�U[Eӕ�&��MUv4��LI�P�c���ί=�ɠrP�~Ykj��Tk-�^��$)�<N�|����ږ����y��JS��m'W�`sZ0����f7a6��Q�6=���Nd�ȇ���Ͽ�>��v�ΣM�p}��3g�#��&�YK����f'O��T��vk�px���x\��VV�2��U���ZYucn���&��6�)&��`��i�+��/6����	�lb9#���z&l��la28YO$��8�\Yf�[�Q�-V��X����(-K��U�bop;Z]�1���P��?ì�cx؈+h��v��X�:�E��e7���&VrY4�.M�y��)�o�X7P���ԩS�?{F�.o��F>��U�$!��+Xy��+j�(��}{�S�ε�miPcX�* 'yXb�!�>��Y��F�,��fNr=�>Zz9~�_�_�`�� �^8��O�^���u�	�S?���BX�4�"h�zrF+�m��l_ Z/�,ō+�R~����=�P� -1E���߯F��W�0V��p-na�\�)�O�S��Do��ݔ���
��(�Vf�:a%%2)����w��i��f��{�&�A�
�n�#�1<6��+�#��'��BV���8�s�]=�Y(�ybB��ϝ;���*333�~���-���ÃQ��ar�Y��*����8�@��mV�0M".o(Ma�!��^|[v��+k�Wqv�C<��f3n��m�.�N�R�,9l�~E�[o���W����|�]���y�NZ-3+kh�:"~/~��L�;'l<��3l�w�n������1��(V� /��4�l�C�cҙ�i��\n�f=��0�,�NO���{y��U�}#{��Yc :D2��ѭI_"�v�Ba�}۷����py��N����w���s��U>�Oa3uX^Xf��#�}�C�F&H��y��Si�Tt�7��-�3iU#w�C��/��/(�����y��c��\Fr�
����?t'��2����吸&=o��Oٶ�Z�W���r��#��+[v�f`tL����&3�Na�T�4��,'���F�T�5jt5-4]���[���y�f�,����?C���؈�re�Օ�|�rÍ��>�S2����B�@]ը���'��z3��mF/�Dg ]j�v�)�j�ҭ7�5=l>��:V~��)+<��3?����$����$��@��f` �M�j�,�.�Hr��B���9qZi�em���\�:���*��:�菄�����G��QK*���Gy�;��҅�,��6Q��t�Y���@#���:�N�V��*��Ⱛ�*�;����D�����$�1���ӛ�ޥN�4��|���u��UZZ;���ه�&��<f� �"]�F�e>G���
>}S�t[IF������n����"�Q�<U ���F�V��d6�H��H��5&g�j���Fhv��ā� �M�>���i�ݪ���Tg{�-��*�4f���U-���PR��OGhGn������G^��,�;�k�ss����|����&��Tj��D�YS!���
�m�ٴ�8[fqA�D?FCo*!���*G"���ݯ}�m����;HΞdm�"C��{��n�%�9�{XZ�c��hj���1k��l���<�Z	�٨���nFߖ�;IͶQ�������$�kK�6�﹝``�5D����g����'pZ�x��l%�ͨ��r2�Y[S��jLn6�V.Q�xY��8w%���aL� �lI9Ď��"�L��ŏ�}�>�C��NN�<���"w�w/C�ʨ!M#�$?KX@a�fg��A�W��T���*�T*e�6�7*�
 ��t��S�^Ưy��A4��'왌�����V�w�tJ1`2 *������74�����[(��P@�0Rr{ٟ'�+Ӆ4y�+vARk��\U.^�o������b�z^@]O�Nx�Z�W��Ѩ��,�fP��� <�r��8�`[>8�"�^Jc���R.��y�>X���%�]��{�P 2�gme�H����l����jVa��m�NL��K�^QQ6�6�ر���G<��_�{qZZ42�ls�}��蠍R>�ͬ���F]uC�����Al�E��1�р�舎L~�u\�N�j��Y�C��L�ƾ[��/�}�/���~כ8x�f*�k�	��4����'�,3�6ǎCw)����O��e�a�+Ŵ�6��՛#\�pY=W^��f�Yk�����x=>&�Vq:��eb�>g�t!&���X�L�u���F-��t殞����B����'��fu%��=���UKx�}�c��[�tu�p$���WXϬ`�����}��\Q���WmA�S�H$��:�2��nm���=���X�A�g�8��c,�>��;ĭG����e�����g��CG�02>���
��q&v�Qc<��E6�ȫ/=����/QW�"�`T��je7i��ft�aFw�O���/��)�[^�����d.�����o�0G���,��ٌ��:�����u��(�k
�C/N/��F�Oů���s�T�K�6�����m����?���۷ށ�k�o3���Qʭ��T	�G���U���$�8�=,67���d�&�s�]��A�6O�����.�$�c������li��Sg`ڷ��=�f���O��ᐖj�F�Y�i���80Z:�j�F+�r]��N�j�z���棐�S-kU�SAZW�1�� �5Il���tȦV1����?V�Ҷ�wK@��L|��BGߠk�Qoi��i�Kt�I�h�W�x�ԚR�*$fC��ڞ�N@a�ZjG�Ag2��x�@�Pea9�:���9]}\w���2
EB3y�
�� �N�]L�<.�j�ZX��ӭ#�]�� �A��S�I�IWnE���˞�����7��:��5����r�߯��uP�0Y̪5@o����(�d2-<�1�f�t	�ՆŬS9T�Ο��}oSZ�rz	���X�L���BSE\iר�b=�'](��	��ش���:C>/�X�+W�[�;%wy�x�6�!���&�z�rM=�g�0����u��:]���%�\�|����r�ͬ%��� �Աе�x<&��W�;�ԛ-R9�u���g��R���윪b����C�x���������رkO>��r�����E�����c��XYYQ���a��J�����(�T7%2	�N���'`N���i��P(L��%J��D�x}
\
P����Y][V��]���)� *��X��|�KȪ�<a�}��Cu�������+W��bZ���gg� �'`R�n�4�Ѩ1�0��-Q"����r* (�����6Z�=w�];��}��/���(�Y� F����X��r|EKg�:�J���֖1%�F��baa���q���h'�P(UU���Wƅ�n>��a��rB{��O�W��e%ع{7�Ϟe��=걝�xI���g~v��}�+�kU������l7p`� ���2�����S����̖�)t�)/��@�b"���T]���*�Qb}U1�}���醏�y�����~�S�y��c�cb�^*�y���yͬ-���/�Fe�Le����o�C._�b�ܳD�^�?B:-,|�ť<{ތ�����p;��5|���niI����nAtp'�����c5&��0yi�r�����ꕟ���Й���V�8@��`qy��s1���=\w���y�G�cmy���$w"R�    IDAT������*-t&3sg�W�$�)�z����?=�_����7�Cbi���3��z�fi��Y���嶷��Ȑ
����>��U��o���?Ʀ�|����z����{Y����Z��fd�N.\�L�U!�5RX�B��kS�;���5�aw*�W��!0��|M�Y�Q��T~�'�#>+��2Z]�J������ｗ���X�y�f#I��Do�P*	9�G�t�9ڭ�����Z����`�I߷�j��ɿ����O���g?�!�N�'��u��g�ҹވU�R����4�!�TQ.`�
��#���b�6>���te�|�J0Pl[��U�s���xF	�\�y�Z#A��Q�o~��t�E�^�&��<��[�Ԧbq�m� m�r>K��Q��d 6�-��k%&a���L�&�I��#4f��Y5��8uh:Y��<���9�Z�N�f%�<-M�bW���A��a3�16�b4ɨh�ZC4�fպ�l6��W�#H��LptZ+�K����4�?~t�=�o���Sm+�vb��tD[�&����?J6�Q���3'S ���;7�H.�HJ�j��B�Q�e����.�Mw{`����迾
X��}��
''��9���
3���^�A���Ԛ���x���6�QU�����huM.�?E��Ǭ3QK�����n���~��~'��B�kiHXk����)��n�{�l�Q*��k9��q�������E���iUh�Ҫk����Y0��b���^���KtJU��mb���K%�hABlW��|�������,��3?A�ZG�Z��+B�|^C�=@*kd=� �l0r��b�Klݶ�o~�+T%��2��<���曏bqTȪ���&M���X����į*�đ-�G@� &�	�Q���U���1���"��Q��!n]��-vLf�O���Z�4)!|���� 5a�n��V�# pp(�+-��0e�"ВQK�U8�� �*���_̞n���J1js&��\G��܇bC��]P�����칰�1�i6YX�-�Ltz�-��P�!�T�V�OaB�}�c'�X iA�H�V�)�}�LH��(�x\N��f��^q�S!���Ζ���*��� �]�1
8�c�ē?U XCax��<�R�����ڗC���g��y�'�r��8�l��ص�ʦa+:M�Q�\����w������1�������<:�e:���K{�:�B�>L���D\����(�I������حA�R0#.qk���3|�o?@(�Bkʫ��m��cqa�rj��Ɂ}����,-Ie;��o�Zׂ��Q��f;ϱ�?����_2��u� +��[vn����s�{itDv`��n��Xy��|�������*/���J>�թ�\��s�[��}��bue��|��]=C���λ���E��Vz���˴uuҕ,����
Fο:�_���q��o��J���N|m;IX��hvq��?���^2���ſǠ��hw�9�w拟�K��� ��ڌ��cht��~y��x�j�Y��9��.&���J!_�lr(�9��Pl��v�Q�
x�!N_|m�@za��A�����}y�￟��Y�z�tr��MSZh2Y&'#�ڮ�)5��n�h0Zu*�]b]�N�b�{#��	�.�|�h�z��A��n!��8z�����j��N�i֊8�eR�W�v2GFݼ�����,��Z�ۼ���s�-��2D��m�/��3<�·He�0���x�fn��ͤ����7��.S��T���P��E�R�c�+3��p�jҔɀ�O��/:F1� �\�떌��jI�Ϻ<Ct��Q��ˮ`1�Y�@����&��$�V�I��u�٦�'J�(F/#&m�z!F8`�P��҈AϨ$P
��@�K�U��Dl%&+F���d��g.��a�yI�~�=��҉�R���\�Z`fz����޻FS���ĩ0��� s�g�P$_X�f�`P�j�7�)Tl���>x��^��ٸ��z��	^�����?�A�<u�j�/�NM�tC4�R� ��#��JRi���
%��dv�
}� K33�#x�&̦&��
���+��y蘴̯/˦��Ŭ��Z�=<D���W_����F��%����� �r���R�:��Q�&<CG�o��|2ùs8��,,N����X@G�é�_����ߍ;����9����c�ưZ�X�V����ڽ�A
E+�6�T�������Z�u��������3=3I���ަL%f�ʹ3$�i5�ת8n��-`D.0!�Rq�Oa����
̝z�U6m���q���
055ӫ���H��Yt�Ō�P��P�O����/�N4~~H�lIi"	E����F�2b������-�b(�%�VX�Xl]պ���y�* p||T�Na{A�:5��&��CO���AU��X�岯�V�cl�ݒL�^�� Qan0�\�1�S��h��-�,�H��Ad%x@�{Hgq&�c���Jz��A����%�P���F��Q���H��G�	�	x=�ՕQ�={S(ǯ�j�툛Z�W�������}���g���c�ŽwL`3��hr؍m������b����
�Ҫ-q��'��c(�����L�^�"zD��F�ʳ�WY ������ԏ����E���ч1�W��ic�Z;��3O�ML)��D��rT%,Ͽ��iⶣwc�;x��gA�$:v Wh�lUCJ�k���$�>�m&�;�������Z;7��F%�F#��ū�_����j��/�c� �쿎|&���'����������/�����cq��z>�ￕ#�ދ�dmm�r#M]S����!5����q׃�ছn���[����sxlml�������شu?K����w���@c�p�����'����+�����,��p�mwnQ'�җ�I-P+-@+C��L���a���\�N�b���\w���!f&g)�T�).]x	m-�C��5)�5ѧ������%b3'�%fiɨ�$!��F�Z��q��+7*MZ�b|7��h�u�c�c�����8�{�����$������&F7m&S.cq��	��&�$X�V���'����!'á�2��*����`�.n��>�.�loȫB�K�*w���T�Uy���p����@r��;���d������9^�\��Ϗ^' +��:M-���R��v���\�4�|�t];C�׮"}$3��Ѣ���Z<�Gt��F���2�R�'���z?�[԰�tJ3�m�h��;z,f����8n���Dx餇]�$5������Bh�d�ܦ�����xu�3�WxÛ�������`�L�p���l�H�(�㴻mR�u�e��>��-\��s�<��t"���d�	(����?��י�_�F��5�¹����Y�:h���y����j����kVvￕc'�(Q���1b�U����͌V��c7bl�����sVʯ��I��c�k�r~���xti���P�����q��k�Ⲵ�4�رu3�RNuK��Ӣ�X(�1�I�L�"�3��N09�/����b%�F/]ÐKeIgs�"���#�@Te��.��/|��=��qy�$*ۮ�����\�3��}},�Vii���>�v�m'�H��8ϻ�wU���f��K/�� Mz�AG�,226�z��b˄a�@ �TX�Ũ	�,{nZٖ0k���j4�oa��2a�zn�^����r�|�`&�/�
��ӻ�	��&'/+-��m��5�{�n5� &�E�c$U�V'O�T�+lݱc�سw��r=�-��#���v\�_e������W]��Z�Ko^e�I��컄����o4�H`-�JbrTPu�}��\V'�lJE����[-��g�e_ϜyU=?c�71?3:=�P�b~d��F�(��A���ty�؋�r�8�ЇX\^�b�)P(��L��?|�a����'>���}lu�{�����k���bַUf����`"���F&X_8���iZ�ynyo�T��l�{���ni��Lry��y����?�Y�����]�Īs�I�ɗR䪫\8�(��"�������L_>���/���C��Gx�癞M0��&�F7�l�r�J��$��c���*Թ]k�c�nb�,�kI&��Xk�.�`ެ4kfmy�9FƇx�Mo�g1q��q
�E.�Ĺ�-��}od��y~��)g�H�ct>�/&��t&�U�:��s�y��	�]	:7cq��F����ɦ���{��@H��������������;�s���sx���§>�J�<�w�Z�2�8�ͷ�������e�{�RL��ȬO�w1jT�^��@3Y����6��$Wh�e�6.\<Eۘ�����D����V�xd�-��c,N1{�Y<�:�n��M���X�U�.$��@��E��a6h�khZMlv7�|\���XO���W���&y���f�΃,��ih������rb^��E��'Y]y��Q7C� �c[8?��S�8Ż��_���mj�6�Z^���Vf�T5��m�^`u���S<�����w1s�
�`0�Skf.��e�S���7�8���� ��8mq�U,�=�s�4����L/��>��.�+	��n�_�G���R^U�G�l��7���~����{F�u�g����r�s7rN#H1��,Q�������Z���0kϱ=;�gf-�׶lYE���L�"E���t�9T��V�}���w����!Q�����>��4��#�n2�������ubi����*SF�a�����?�x�K���ES&�rV�iN_����`ja� ����bY�g��,>��ql�4�V!׿���_�dr�����F�o��j�ϭ��~�5����}�)j�Ξ��z����y����� �������G���O�,^�ŏ�k���"|�������?N����M1Y�X��P��s�F�l�����ij�E�.�z�� S�@�3Stwt�Aa+�FzE��I�D��H�-�UEv5����^G��#8���YA��UuܒGW��2X���}�D�w�ѧ���"����@��T	m6�� �F*M�l���(]��������F�U&���t���F���$����lc��4��s3���p��;'x����[[Wc����v����چ�u�Ţ ��;y�
�5�H~8Fm��Wbj@-�-�P�mFM�+@O�����x�&�P����uI'� 3a���0}�a��^Y��pX�ܹ[��ɴ� 
(���E,�\a�5܌�mb(Q��D�k(`M�ۦD�]@��~��d�&# ��vsll��2����*̧oV�	��)�	k�����Y�D����.@R^o���
������Y<.�b�e�\Е��H6�S�#x�{�U����dhq��&�gN8��������;os��9�6{���y�j|�����*�s��������3)���)��k�ְ2���w�e��)�g�qФ3⦳�C)� �q���N�>O�`����w���z�`����۷�iq���4�M��&������Y����ǣ�>Io�N��k�ų�1�;JW�n�V��+�r��_�d�nh斁^��t|����p��y����q���g�%'����J����g��Ͳ�4���4����w;�<�0T���O�d&U�����>����tl�o�͟�,-��ݥ�O���Fl�ˮz�� �ʧ�� KH~��X�/�x�G����%F/w=�{������D9*��?�;�����F2�;4���5��{�#8},��8{�>p7��*�N�a�VL��H�lH�
�ToR���;ĥ�y:��s��Xm:��2K��=54��h��<����N�X�_�P�M��P��z1��mU�ڍ�N_�z˄��χ�(<����pq!�SO=����Cwcw�X��`��ìǲJ�+�DY��Vc~�$��8#C^%u���Z���Ͼ��<���՚�D2���v@7U�u�� �����78s��}vl��<���)��S�5ebH�j���])�:ԃ\S<4�R���Xqw�X5Ӫ�0�+�Xwn�F3��q�  �ז�#�YB�l�jJ+��-�؅��ġ�,OMbj���+����W����Z!�_W�k^s�J�J�\��I��Q]?�40�\A+�E<_ara���
U}C�h�<J���_e׾�8p�fܞ0���d����Q��:N����O\��>�n�I��dl���3��d0X��<o���j�����u����(����kK���G�����[��ӟ��y=f�E�j5�FL�z�G�h5:{{P���;b���ŏ����Ǚ�/��X�RH'qh5t{�jt(�a�O��j��6��u���V�D��d[t��qvn���%B�v�a�e�[jhqaf�;�Xn<�*$rmݣ����J�T�u�y��GCr�9b�8���&��(����=�kBQ�F���A�����ǝ�*��<�T�F�J�Y�k�>�'x�[?��9x�~v#닳���k�~�W�.S���W XCժIe�*��lj��f�������uw��|���!n�_���d�Q,�� ;Y^Fg=�]J�&��x2�����Z�\�
L���G<z�(�����8�zd��O}�ӧO����n�P@�6���U�%��S�+��U �,#�Q�ݻw+�ťK�w/ n�/[�!�Kҿ,#���C����~�>�VQ�R�� �W_}E�_�Q���K/��!!�
�#�h��'K��:C��ψ���O��@�L:����{L��׏��4��-9��+�j{��j��-ZW�JG$�F呀�_��
SW.����b׮]�z�u���XF���C��/��4��oU�����tw{���E�.5Z2�"wP�$3�5�:����d����2؉V�Q�U�Ztb�]ݣ$�f�����1˫I.^�B��b���R����*�~�ݿ�QJ�s�^~�w����WοN�4���Gn�<��V���_���O�u��\�Y�6;��N�������4O<���I��7�b��V��-��奫�5��S�c��y�����n�ZH3{�]V�^g~i�����{3�|F5v,L�$���pu)�=_L������T�>�|�PgX��T����c�a�Ь&"=�$FS���-��l=L>�������f^��	0��n���]=�w���n���5�̾�7*�o������'"�6M#g�+Djc��ϧ�)��V��f���
Go{��O\�ϼ��>�Yh���>��^g-9��W'�)p��Gx���/��Ջ���8�� m2���Q�%UƧ���z̀���٬�u���}=�;���p��z]�Ё���l�ku\�2�x�\'�t�l<���%��	:�&L-I;�Qo�xy�-;o���F�B�6�ӪW�F���O�S����iVVƱ���}.���Z�,ּJx��+F�Kذ�S��-`�kؼ6r�"�\	��������1��z�@4�#���'9p�:j��Kd�g	x�8�:��:��E�P�ٷ�+L���ij傺���F�����8Kfy_��#*f�&�����@��ʢ-�_	�6�4�k��%��<�n��R��}��i�\����-���Q�iM3�bҍ*����q����X]�Ȯ=C��&��^�Vݠe^Q�La��e{3�{�W�6��5Px�}�3�@������/�짅��>��T�D.�"��c�z���F���-j������rY6��(�V��W9u�5F���;�Zl�URuV�i��u����+	<~z���;z�Q�va���(>�4A�\!��nl�w(J��VO��t���^e�-����"�^���=T(!�¯�15����h�����T�_�!�ZnT=�D
�jV�k7Ŵ���5�E�u�J:��p�{�U���F�?�6��Zl��_��b�f�$�Y�;E��utu*�N�k���S�?�EV����	x���d��]����X�- FF��Љ�/
+2ue�+S�*�F:�7���m��N�t	��e
&�L�ߖx�'�P �֭[9s�̇����yM�� S�٬�S웬['2*�ʦ1�lj:�i����ʶ��)�O�]����)�m�kL!�    IDATő-�)`W�$4W�+�L)�%�P-zE���e<-7]��� #`Rι��ĵ,ൻ��!T��������qÑê�����_���z��J�X,��&O(��[o�áY[Y�W_b׮Q��E�����2������*^T��Tc���R�ӪV��,-O㵛���R����"�(�$��ֻ��������[�202�j�U3�J��p��9���X�����r����`q�e�ǟ�e��0�g�-�f}e��_<έ��@� ˋ�"8�&�E~�ӿ�ԥx�3_����������o�	)9�8M���j&FEOQ���-��؃|��Gɥ�\9�.]Fi���/r�_�n0�[�P/��ć,,�?��L�BJ�Y�J�*1;-͈��Q�Q��O�!#@��=4�:=]a<�u�OM�+�������>I�f��{��}G���̏��F���7��䒰������嗎36�Oo�K3��k~��Z����4����L�R!W)�蛍|����!b4�!'��U��
��Z
�be[�<t���ߧ�E�j5��Ԝi�k(�6��Sƚ�TJ#�4�@"����b��<�3��j��'��-�{�P�F6���u-`&=���8���$�qhM�;u����;�7�UE�(�^�X��i�{���2�\���9l��;����kص4�Z�FˀCsbҥ��J�^o��reU�(��o�a�<��?�����i�Hfc�tC��фfw`64���E,¾�]j���ȣyڕ�ݡn�����)lh`�;Yϖ��Z52�U�������SX2�����)��H4Y�B�ܕYU�����*&��JJC�hh�m��H��v���*V�t�����Os��I'ױ[���:+�1�J�BW�[�;��!�a����C[��=����
��-��@�����/�z�������n��(�r.R������b�y�J�j&�*R-׹r�<=>6�/che����nw�uhŊ�[�M��u6=&\]9�=�W�Q���?�h��R���Z��<5����pݎ^��uu#��A�^hb�J[C�\�](.;�IXBi�(�q�����&��&��|�@�+:k��J�&a�*��G�^{�/��&�F�P L)���G ��P�.� o��r>ɛ��J��2�ͪ�2���
4K�V.���\T]n�%�
`��:��$$U���չ���	�v��!�?��/`H���r���R�V��d#W�h˖-j�ܮ׳�_�J�S@��x�q�tK�����F+�AZ^��p%�#���%F�%���R4��8Eo({�A
ؔ1��QV� b��+ݤ�Op���  Z�/�T*������cw�8
�L�S
�8pH�/�Ѳ,�����)�)��8�w'#p�y����=e�-��?�͡F�S3sD�!�����lVƟ￫���p����z�|^�;���*~%�{��ю ��S�>lVхԨ\�.g�믻w$@��ar�r�KOr(���3���ϳ}{7��*��*n���%9�g?���u>8{N1V�`�fբ�Z;zy덟��+?�_瑇>��x�bz����I��������x�obei�{�g<�ؗqy#��ڌf�7��?��7�4}����;#�;��_"��c��	�ʦ�T��v�^x��)I�[�x�O>�9��1sgn���1Gs�O����l��X�YCo6p��}�@�$��-��'�Og��e4���Ԣ���|<O$���Q+�07�$�O�P��8��q��'4��s:�|�Oؾ�z�&��G?��Wf���?F�bc�?������}L�	yl��Yj�&n��t.�4n�J�l���#:2;ao�x�3�����������}#�����D~��&���̨�d1��iS��|����bm=N�,�K���n+K3twFh����[g'��X<���ʽ�|�;�z�l����@�Y�k-���`Mf���g��dr�ˠ�Z5��BNz�w�g�A�ݓ���U*ej���"��P�b�[��Ģ��ٿ�Or\�͖�l4k-�� �q*�?Kⴙ��7��iv�W[�E�g�p��F�A���Ⱀ�U(��6�F��ˆ�b �J����zzF�)�I����hTSjk��(6[$u�\{q7��DS��f�c��*Y�͆�*�{��h��DB��ψ�1��������gt�� �D��>����C��/���4������x,�y.��r.E#�Υ��WssI<�*e�26{U��̶�Fg����e���k�����gࣁ�3��p晟�k{�%�(�Jj��Uٶ�(�@'������>f&E.��*.�/��U=F_7M��l�����R
w@����)z;�x\M��.���EK��/a���4�,U��ń���;��R�M�k�Z�jK���Fq�5���!Ej��jE���EF���XMe	�2٨��+����Y��~��*6W�������_��L��y���? U((P5�׃�nd����K�gd?]=��w��(�3�bY)�ج@��z��}
lT���t�nj�6��D�&a��z���͎ ��v*�%6AN�8�F����>��ǉ�#��CF��	�P>S;�ehHz|�! FFڲ�\�e=���r�d�e�����+�P^۬��O�% M�!�-`N ���
�yEXD�˘U�� e�d��0�r\��$� ����C�
��ݫ�P�en�2�zE�wٞ��P*��x�FQX�����.Kj�D�(��n�G�Ȃ� �C�
(O\�T#no��ŋ����19>�O|���E^|�E9��9ua���+�V������*�����]���tYT���b;vhlXbC��w�ʺKRKY���/�ڱ��aF�z)�Wy��@�1G0b�Xob6��9w�/��\�W^{�c�|�b���$9�U�y�/�ũ�ߧ;���t�/�6��N�}�;�b$����0���L/,����[�=�G؈���7�jI�|�i�!۵o;�_��L����Ųj����banV}?�v����v��Fy��'�kμ��|5���}�,��o��׏;�k�H�cX����z��7HCth�]���V;&a�R3�#�M��U�=�*	��X��i��p�4��4���ԌN��������H���s�͂b������:��k>^,a��Z�bA��F�=�9�8mN�^��!&�t�D� N��͍�a#���ҕ��!jh� W�.�u�{_�3�^/gJ�������'�Y���P���w��,��S�/y@X_�bۖ>����ίl(���f����(����-�ɗu�"��Z�]5) O4���4?��ߒ�_��h�O��j�av)C��-[��V9}c�K�� ����aj�W/�2�ٱ���[{H�L��h���F�PE3HD�+���I<+fk����,6�jI)�U�e=��f�Ҭ�9]꼈F�#�UN^�u�B�%*�ma:;��+��.c6Tp�J��:�B_W�ޭ��,P\^�'�EsJ�]E��0+���Y��h�[6E:������#���Õ�	��V�<x�[��.[q���Y���]]������$��N"gd�
	^~�Y�C���� �������������݇v���𘄈^��v��gࣁ��Ϟ��O��Ԟ����,-�L\��cw|�ͣ�6۶D3GH����4C!?O�������Ξ#G��:G�\�e(�|��dm5�>H�k#��aw{T�c���/����2��)Oe��o�����IM\U�-�ֶ���Ĥ�(��U�FR�f��<M����ѡIՖ�xn�,��;��`b���$��6-܎ax�sX�v�{�
Y#Ǐ�G��G�OT2	�Ɏ���&�o�~����YK���&%�.�Z¸�,f�l�#V@� >%���1��H���-���:{��&���_���a��/�[��N�8����A�Pk�(��J�&"vY�,#�Nb*��v� Y��heD-�+�X@�&� �{�R�*&�	�V(�����䦰���L~d$#�/ۓ��(x3�P�#�a ��]�Mx�T�C �n:�RUq��v��䊆s�#Z�!d{jU�`�Pc���kyO�,暄r�
��D;��ۥ���gaLʅ,[��)m֙��T?���J���)���L:�Q��_����6���O���?L��Wn���	f&���'�Ui��e�|��M���������m[سc_����~���M��A����\���w��'����"3����'U���jS7�tq�^�W�z�_�H]N�?r3;��1��|�l*M��C��˫o�ͳ?�5���>�3R:�p0�Ő�{���\�H(lR}�E=@��^��=�����8.�G�T�:{�y�����U!��E�fh-�����Ŭ�_���bMF|V����ܭ��DbR�3����*�{�!�� �@�:�_���^m���Y[Y�&�z�F���P�a㙭	�������*7��Z=�/��s'_�VM�u�#��U3�d���F�����Yl}�D�4����n�P���t�Pl�(T�*�����-�Ē�4���g���{x���8��&/����L9��POH�rـ�`i�@:_&�P0��<��[�7MV��y��WUv��Z���X
���p�Ǖ�9��1Z\X���$�9�������:gμ��*u�N�l��><��)U�%��"mA�����f�Ti���%W'��r�����>?��i�^/^���ʢ�(��c�#W3y\3���[��j���T�ʈ:�\+�k�|�Dߛ�eս�e7S���}$s�B��t�׻���J�Qci~�fy����dg H�TS.s"��*��4����
�IK�82."�ѤQ�b0���@�lQLfK�0)�
��:7��m7rñO���Ӓ�����e#S.*�U)^ ��b�j.�樖78�}���L��'ґ�T^Q ��l9<�z���k�4�n,tm���G�ss��O���O���I�cXm>֖�>3��=Gq�"�M��8Lw�o��.�\�J!��4VkU55T�E\a�W1�y���T%_S�e!���ׄ^+bs:0Z�����v�(t&W6�{�حZz���L��<�Z2��m4��D�d���U�4�T�l�,�"L���y���	�٤�ts��8��D���ZᦣOp�]��7��k���ɦk�<u�b���n������2�} �jfk�65�|��������G.Z�����G�D�'q&2b���S7{x��{��J�"�P��ͬ�c�s�=�b����L~�)��ŕ�V\�媘bj
<mIW
�&,�r&��	�&cX�0' KZTd?�ɿ���7�=�aی\{d,Q6}�jYa����dy���	���;*�A޳�}(�����²	8�*�u�M�',� 9Y^�Go�e��l�\�Fsb@@-7za,e|&ۓc�}غu[{�	����o�ã#j�\�0�&��)�B\��vl۪�Ybi,�
���c��������4ӳ�tuw�/��M�m�Q�믾�}�=���,�s�;；Hg������~�~�i�x�-����\|���k�=��S/2��geq���[���p��8V���}�h5LD�H��|�_g��+�ty���%�L�{�~�n�ce�j�H�;�9Ŀ}�yVV�y맸��G18ݴ,&�������{,L�ɱ����L�����VwH�+�6�.L��o�QLI������J�]!M��� �����E����b�+�/��	����щ�H���\:E�\������妿���2��k��5��%��eJ�,��� +K�J;���{�>��F�륜MR/�8u�M._�H:�$�o�t�Z��?���[�ri��z���h���Na��5���ɮ��YZZ@�ٷ�4^_�[��I80�����c`�7��'�"e,�4ֺ�V݈�⦊���K,�W��l*�h_T1��[������#�#��Ӡ�j���\�Ǳ�ݤ�:NW�jʐ��V���g���S����q�&sK1����⎛)Q��1k.Š*`�K��Q��n����6Aݒ������.L�"n���Ļ�®���Us�n�(m3�t7�e��.�9H,����C�\U������CK^�o��Ⰹ�X�V/a��
�6j� f�����
���Wp9P��M���d��3�O7��u#�X`����c�U��4�m����P)%�LVb��F�r5��3@�w�rJOL�a��y��/�,U'���ޠ��F*��P1�X�Z�@���QX"���ʌ:�r��t�=�9�U�$4R�8�}w���c���!�kgࣞ��
W�^�p�;?�&��b�)�Y�h��sX-A�{��w1:�#v^�嫪v-�s��/ ��Z-��o���ilNC}�LON1:�G:��Ԅ��.�N�QBs�1k
������re-���P���b�K��!��J�b�n�Ӫ�h�vJS�I	��j1h���KYNE�'B�l�7btژXXbb#MM���{ؽ��;��%B~f�,�;_�*��%���<��}�{��%�����.OOc�Y	�����᰹�Z$�fE1R���UA12��l��d�6Ú4ڻ_�%ES(��nS�V���B�;���C��T���^%37?�4�G�Q:@�����C�#�%?rCp%��0�� �ݺ����6$	0%� �# L���K�G�!`H��a1%Q�����#73�ק�_��	���"�ݙ�:�F��h����J9������)c]ײ.	��_*�V̄ E�o�x��0|[�#�S^���SуʘW2	e��RY��@8���j��[]Qc���^�_iQ��G�\Q�W�8[5;�R���U>8}Fu<�k_��[��s�����.������ԉS�!n��c\��"K��R���eum���s_x��{�|�����i�~-��{����u�j����nf�̳ud�J9������7Y_<Ϟ����:w����[U��H�l<��1[�\�F��h0b�[�H{y���]�2��F��\���i����W���n��W�x���,9���}DzG8}�=�륧����������i�m�eUƐj-�$#��_@���P�!��6Y-��555��X,>崕�?����)tIJ�,MS�"���h6�(u�63��YW���*(�N��evvF�3���L���:�.V�Nci������+�O��t�4K��G���L�IŬz����K��B���&8��+��Sϰw���ς�-��4�:z�q�l�V��47O4��ڬ�:�p�N\��(5}4�N�}�m�{��WΩv�ox��;��:>�C1yնs���"�Y_��;��:��ƖdӖ�YH��c]C\��:*�
V�K�kZo����Ab%6���3h�!���Ae�����)�z@ϐ�%�wt���A�|�ID�uժ��ޤi0�y(��,�=����(��N��*�r���%���J�L�։7����U�-���}8�-N�z�ׅ�f!S���`͖(&6�xE7-]�톢RӠ21��v�I���iQ�����L�N�v�i����|V�w�H�oYqA�m�JE,B~�,��{c}��� ����J}��g����ɔ�ټ��SWW�����{�r�����Gז�v>(���Aߕ���D/����ͬ�n`4I$���f�M��g�h�T�8{V�yLj(�m������rM՘aA��j��'>����0n�D6���e�.�_���0C�.�������B/{��b-/�QT�X6��Z�A��2u���紣r*��wbV�T�S�&ul3~��=F��T���Z������w��J1������ȅ�����/��.�K��������@4� ������	֥ު\Q#m2�lw����
`��L���W�b���7ݚF�$3
��ڶ���~�����y���Q M.�b�P5x��͓H12��L��9�
P	�Vj��XF��8
`��5r��)�Q��B�	���٦6Rn�G ]۸��   Q�vrh��#@KΣ�u��4�~y�����0��!��$�Z���B9��q�'ˈaG�I���_ar��r)p��V�	%�$K����%9E    IDAT܈7�X9.�:;���fs�/��R��Xm�ƾ��� �0Tc[FU�z<����(��J<�T�W�xGF���F"um��'�K���G��^5������򲺲�s?x^��ʦ
����gy����,p��::<�~�>8�"?����l��c����_fna��L�\�C}*��7�c��v�HLb��y��c�d1�1����:�����'p����؊�&���y�X�FVg.���صժ��O].:L��������*�r�r1No��ݘ�$��f��,�ͳ>u���{�؝O���T�������*���baa�\.����{�z\��>���{;�D(�ZL~4k����4J+��B�����z�|����#e��CI,l�._��L:�`nPi�I��lĖ�
i�5��if��H�׉��i5����p�qw�THPC��Ji4����?R�z{�(��:��c�B!3��W#���R�o�Qʗp�܌lߍ7܉��$OR/I��Skj�P�E��r���Z�:˳O���K*���c���論F�nR��hG��+TC�0}�~����ӯ�;�A�l�(�ghG��Vh?`Y��*�Y��h�(�X���	��&��>�E��S�]�*���ۥ�誮����Hg�tR��)62J�Q-�1���*Z&N�K�m�z%�(�z��o�ѽ�2���]~���b椽��������%�<��۩F�\�T.��C��-���R�R��@7��UTI�����¨P�ЛJ���+�KM�nj&;��h	0;�F02�m���E�0V��Hƣ��@:�F0jgu�
nK�V#���8�L����l��՘�T^��Sk��}w�֎�oנ͵3�Q��G�33?�|�;?.g�8աk4K����d�LΠ��;:{w����)���<�j���Q��g��;�+=�����j'��`j5���cn%UՑ�-L�z���f��E*Sb�Ta-�!�O��b4)���Ն�i�%�Rc��ʽ��Q���%�/���D�{0Y�	�F��K�˪6N\ȗ��1�^�j��O�'�z��'�T��aadl���9~��+�-�eٽ��~�#�C��/��k��	$����x���ۥ@��S���7�� G���P΄]��ɤ�,�,��Z�w��R� ��`��\^���|���K푪�H�P*�� J
��j��,���#@IX4�\lk��jY��o�<����/�G�E�}��+Ea#�˺�G�]�|�% �X<	['�NΙ����1������	 ج����s,�,�T�#7t�
�mTkd3鶓Y�N�佲�p0�qU]u��������E^�#
��/.* .�c�z:�\�t��hD�˷�y[�J���#���2�k��d*ù��H�3��,=�݊��s'n�����ڟ�?���Y޽w4-t	�:x�g�gznR=tl�>#��;k\��+��*�b۞}��0�S��!#cc��y�C;n�Բ�0������9.\z��B���;��ѬP��a4X)4;�^�9qe�B�Ewp �7@�^�t�L���N�Qؘ��G |�i�Z��1l�B���w����?��4W'O�ѽu/�.OQX���s_�C0������ϱZHsu}�rQX�,�sW���Tz/� ״�2|����d���9D� ��ηX�{��E!.c�u���c��/�YTs���"�/����^��Nb�90�̊qnU+4�M�M��4V��\R�\�w'N�������OhxY����ۿ��_S�<�[�|e��C8$�Z�`(R��U�,o1H׭dTT ��aUL�hkMV;�]O�l�T(�z(��lm�wrb�ل�g��G�������Ϟ%��Qkp����{ϧ1�\��Y�f�Ո�ZW���p���q��oI&uUՈ�"R�W&��b[�6n�w=����0��u	���J�k�ؐ'II��r�ti��ۺ8�-J&�@�)�>UרW�����J�\�Ro��V����1Y,���}4�Q��~�O	�bN�UZ<>�j�&7H���۔�?�̠�̸���lѶte�Elm^����8��|�ݍ�i �<����~�'Uvi���aը5�A���<��i&y�7Si�ru�B̀�!�k2��&���q��9|�.��atݬ"rlv�BE]+��.�������QO���S�@�����9��8{�b���;���n�p���w�1�][N��G�+3?�p��3�9�u�y�[���@t1X�A���s�tJ{E���ܮP�Ӷ�+F(��"�H�	��6Kߠ�Z#GwG�AG3�1PU��u��-0���p J6_���Uќ��t�t8kx�&�|�&o+u�����0JÃ�VJ���Uڼ�и�U��|���Q��������>�Z��ȶ;�����ߟ�w�Ӑ�mÌ��ƫ�����"'�j��=<���A�2��j�2�t�B6� �tBˏ�$#Pƭ2�M�c
�u�H�[[�&���E4����^Ղ1<���W_cl�t�y��ߌ_�������%�pthX�lJ�v�q2�V�	�����@�����v%��A����R���ٳ
��AE^�K���G�����D�P���u\.�d�ή(���D�C�� �M���K�Qz�g(ۑ��{p
S( W^�Fm��BY���e��-a$�}E@�s����U�Gale���v76�j}� #L��#�|��P �l_~����W�~_P�i�S������|>.���a�x��x�����O�����nQ7.	+�y��)�j��ٍ���{�S���g>Pl���e�N�|��-#L/LrӍ�qp��j|v~�,�t�j�Bbc��n��.�Au�ӳ���/�/<��_��^�e�y����н�CM*�.��S�O�ܥ�U���l��C7r�h�WU�rt�NM����If��3���$W�cs����6�c�'HGH'_ʱ�� ���{e�H0�ef~	�iS�`��FSO�D���\����ȱed=��HM��{�()�#B���2��p�rWku�����sԪ�,�/�O~����$�+5�|�M.]x�:���ڳ��h'�m=6#��^!�L`��qy�*� �M��+E�nV����n&��#���Sﰱt����1�I"�8�CV��>��'y湧�
��V8tݭTjF���XO��λ/22�Z�`1��E#�\U�E���v���IY���7��a~fs�@�i�/����Ru�D�������*K���ש��hf'�{�뮿�ťu:�Ĕ&Z�
&�n$�2�y�~�o��:I(�B��*�Y �h�v����0��8(VҘ�5hT�)�ٮ�|�b�˓g��l�e����V�ky(+덶�����}~��<֖����RW��Z�E<���`��0�Ta!�A8��&�����Ӌi�:�n�zU�U�*-�w�҅�+I,��},�etc�9ȋ���W��5=G�nB�	KMg�@�j�)N��Q�Na�*�(z�f
z��Wf�wvR3x��4��>��K�t�pG?��r/6g�X�栘˪�Q�'��>Lr~�7^z�����sl$�ٳ?
ʹ��uF;�T�SH�1�'�x��z�\;�|$P81!F����g�K���v?��\�L�ӽ�����%��Ra����W�Vh����i��ಃ���b��ta6I���N�%͚Si�Z�<��Q�A�%��s�	�#D<6:],ڤZ.�s����!�RUZ��z�n�!q4&3庑+3+�|*3��߫��p:
��q�d��mw|�{g-�bt�*�*ހ�W_y�ŕe�s:4��ʡ��SO����*�a��*nP�P(#T1jH��0fm�Ѥ��*��T��;wN1[r<�dV�>q)�ŠV-����(zIY� ;�#�R�/ D��4NH��6�!�R����Ü?�7�U���.̔D����^Y�&�',� @a$Š!�l_�̻\��������0u�#i9��T/�<96����6;��h"�.l�<�8���m�
Ж��)`���[��7G�4e�*Q;m�rY-���"��4��_D �c����;WP,���`^�ϊO���ڊ�P����~q��lR&�}I|n��tuD���9q��;@�{���JY(��¡Sd��H���-����T�cǎ�VqMOL\�g���ϼ�@��ݭK�Uf�g��tb�H؇����!;{vtP�ڶ��S1����
K�s���nW.ҙ�	
�ɢ���8=N�?��p+��:��
�D�ޱ���㟿�}��n�2�!2�N-S.��Mԋ��D�2�����4��+܅'���*`>4�S}v�۷�Y���6"[���7�eme����}�g���\z�u�n��������P�m� ��s�"u��x�$~�C3FC/`4z��cc�y�70;�J��5�y���Ґ�b���榮`�WH�o`�l* ]:�+r��p���.n��T�Ŏ^j���PA�KK�<��?PJ����.��,o��9Lh`7������b0�UR�Gj�8,F�[0Z
T�k��΋�]6՞���C2���kRM'�[�"�t���#D"���2bN1}�=ұ�u��5�ĝĉ���K��U���ٟ�	Ѱ��l疛�����DȤ�8].�z%�î��2ų����0�E�ml�ϔ�;v���Ѭ��f�Jq�]��m��|�
�>�����Q�W9�o�����,�YZ9�Tj-U)��h��-yv��֜�jR�uu��jJ;���I_�&��$y 6��E�
�BQV��
Om�a5Y��,'�}��f�MS2�x:O���0��hVU���:�e�~�ʺ��ue����hb¦�[HÒhU��U�Fy��IJ�&��1旊x����ʕ�y�m=�7}�\����[�R+�K����Krkqv����2��Cߠ�bq�A�nu�zI��kY{�v����\[���H�����\~�G����j%�t'���9��J���f�R��/�_���j_�b6��Z2�D�����h���X����P� a�eQ8��2({����1������9	k:��j	+�Z��rڨW3X�q�c����Fͧa���TA�Lv��N:�J,'�o���be%��֛�X�q��r��>|��eym���
o���Ғ\�������c�<D���b���T�K�a�R�~��6�4r�4�p@]��_��<J�����<�9ϕ5d̓J�R�$UY�%Y�gam���~<����0�Ech�q��xĲ�eْ%YrI*U���j�*�)2#"c���9�T���V�U+�"�������>g�-�� CC�	��򸕑s��:�e��|m�*�����;��jQ����z]A��~��y]�ŋǫ��<��}`�O��k�rf��+���Fԙ�
�:wa���IZXJ�NƦ����Ty��[a��a#�|e���1uv8�����RF0k�$�RIA�C'�J^+�&R�)�$�+h�s  T��އ�F�����
r�8}}�
��;����PƼ���ۇ�a=��:??�`w�vN �(���n�T�S�f�;l��(��u�f��KW��X��4[�L�lZ��z�N�>�ŋ㡇"���nI�Ү=���_�����R5�Ip��9�����f��=�w�]^�u<�C�;��*w�f��e�&G�� ����?�/�S��g�+҃�v�)��<����K3`?�У�`���%��n�Tؿ�뿆J����������Ȫ���&M*f�پm+f�����:�bKKo��M�e�	{=�u3�Z���A�.z'���ǟd9��3�Ǉ>����!ξ�"��u�;��	��J��#�+������1�^��u,�eى�8L�`���fq�tmQ=��l%2�ǅ�o�?��,��`6�uXab�v��7��C��'��lRխ��}�[�i�@�/���ص���a��<~���j�Cw�\�ύ�S3�$�3�v��~~�?���ɘ,9�^:At�
{�nbma	�Ѭs��i�Zo �z)O��`p�6{������~�k_��[���G��(w�<�~��o�-�|�[�����b�����[oW��f��i1J�g��H���,����|a��:=t�Kq{v���w���f��M4�],�EWѲ���B%�J"v�Z���	z�OvMZd�����.VIF���Yd�����ڲ]��|+k���{����2z��������8�\~��@ �҄��0��~�V��:����`�PF���%e�����-U�-'�9�N��a`,��&�o��:WH&k�b#S*)��9����Ւ��jJ�E�N�#�ڕ�u;w�n6���iT,-M�Ȭ�cD5U`~�&;���@�p�ˠ*�j���_����������������{g�ݞ�w
������}���K�8%��P�޼R�E6_�ɠX��0���l��hӶT�[M�Fk�j��]�V\�6uC��h�|�4�-���f��E��������\�\�Eod���A�����S���e������JiH�I���C�!�1S�	&v��gHՉ�B���ej��L��kK��v�F2٦���m�FU�R9�~M�8s�e��?}�p���/���w5�A�r���L޼I��8�xR��0@�ͥe�T����,��6m�T��ltL������^�5���gMb�d?�8	�%��!,(��'���w��6
���!l�F��l#�a��+�P�]$ܭ��͵c(��� %��D.��'��F*��[̝7�
e<*,�$Y\��D9'����/��l�$���5�m{yK��R�A�}a!����fM&r��(�[*uƟ�
{$��Ҷ�l/f�2ƪ��u�I������.`Y��ڵ����Nߔ�f2�&4��F���'9t�A��y���Y=���ݜy�fS�e�-%_�SA��0
�.,�|v#cc��y��E],��>�[�m����'��K�Rm�y����	��Gj�<�O|��nM��]�a�l��ΰ|��k�qz���+�s�u�:�Ipwo���Gؽk��{�'d�7;
�� w��qej�旸t�<�3�	9�l	Ҭ�)��mV���r
�ͪ�#���?��|L����>2�����.j������ę7�[�bp���``?���p���y����,�0�;�2-1��(��8�V�� �����V[���h��X�Yxm6J�k� �]��#��eL.;W'/��_�;����G?��\������_���j��C��o���9��in��v~�ӿ��i���,���ab4L����~]��>���\�*:9wi������
�>n��N���13�R�R˸��&3�rQM��~ɉo�.���:�bb�Σ���DW��Ww��ˬ�L�����Pz�a�>��m�I������}��
��Ç �fyu�'D�+���,.�U��^}�˗Or���f���x�^��?��`�^~�8z�n�X�6hU�(1�`tq��I��ij�$WO16����_av�e,���ŋI�+�==Ԥ�ܨaŌ�b����,K�>���E:[�i2P���璄"A2�V������{��V�E,����\�B�fd��{�_\e��e�z���NĖp:��9��a�ڤ!e{��\+��8TL
��s��������Lb5cf-��{B�P���
�����R�������_X��{_0���kl�6F5��lnP��Uݽ<3���f�-�(U�4�I,�:��X�Y1��M���{����x�����;�
^�����_��˙�=�~ҙ����|���awS�2��[�����L�M}u-��D�ͫ���&��l&3n��b5��fRT�Ѡ�I񃳺|�h����lbkh@٤S�1�=؍uF�6��+P�Q�D�8�rU�SӡB��m{XZ��q:��=�,�av:Y��2�Ej����^n�le%^�l�`��՟p�����Mr�y��y�z��1��o�����b$�3*��wOeu����	�דx].zz����� A@���`��XRo4�<Vo�yk	�����1��X��t�W�FCK�"p؈�P(�)�H�]T�ew��X�[' K�3�=Ob_!���F�Q�&�_I�&�%*    IDAT��A�.�/�
X������5�_a��i���~ǴZ���;y��]��q�sr×��x�k���9�(���u�\Sp���j���HCK���%k���U *^l�� 6�*��(���U�
"3���F�s0�W�����������ul[]����s��9>��Ä�A^=uF�10<D2�cf6���ū}�1�niaQU�w�y���=^E�(F��B�d�ä��M�K���/�D<�"�ӭl�7��el��g�N�)���[���J��A*�n-;Y��,\��Y"��6��bdj����;x+�B
��^�1~o�������ŝ���G=/]���]g��O=����e.jR���UzC^�,C���r;��^څ<��2N>I5���X��1�ݽ��_�(���n�У��w� �����gϞ`׮}�u�8�R�іd��^'�	I,���N��-�I�gh�L_�0.f��v0~�Q��9v�Փ4J>�k��^�������gia�?��?d9�DW$��e���ٹ5R�}C�j$���>!��_��c�ط��<�mL�~���Y�v����8zx��d&�P5x�:�����y�
�����Rf,�_�j�����M����:[$	��"�`0x�W�l��.�F3�s�
�׹6y�C̣Ť_l��Z(���~������O�|�b��}�|��s��U|���Q�W�9�D�V�N">O<1�/<���0���SK��'�⡇�����;��-O�t�	ur�o�
_
�I��i"�e"� �|���(��.���*��6>,�K��S�y�ND�_���ئ��R���7@��������|�N��[�]�6��Z��U��v�h4�`��+��@wd'Œ���Y�>طؾ�WS�҅��V�� 驛�\�n��d��I�4Mb��l���	��	5ZU*�f��B����e%�dfi���b�_cq)A��]���cg�N���f�>?7n\d�p7##=�~���4%�V#�Q�h���5��[s������A�����=�
�^����S_��l����� �\�cm��ʦ���f%����-M���*�d�%��r��jcL]i����ܺh֚M\(ޮc�֩5�Y�Z��`���l�*C���s�����|ԋY&���lc��em��(�o���>B=[iTژ}~��<�%E�A�Y�*�U�M��=���x�ko���j|����mL�+�.'ٳ�v�$ׯ]��Wk�b>�ޭc|��f��[U� Y���^�.��͡@FJ��}�d2Y�o�o�rQ0�!��jc6R�H���f�2�M��pz��$��MO
ļU7���)�Q�N-��2Y-��L��ZZ=I#�.+^a��y��O%�[l������pXA��F��C>GI��N�\B
�l���gU@��166��'
�,aa
e�r['�QDBwg�)�Y���-���l;,�7g��Sq���\N�%�/�.u��$vND�`[^����DX[��\QA������s0�QB��u;�9\.U2�+�(�'�(�E�����b�\S��O|�c��9Μy��߶m;o��D�พ�z����V�y��k�|�_����\�@8܍��ӅЉ/��VT�j��C�J�\c%� ��S��$2�>�}|�4[��,��r��g����	�+��E�0��t�I�M�r����*�L�j��g�sԋ9l�2�^%��&�s��u��A��;�z�A���z���Q��lⵕ8�ғ�-%5�nU���>ɜ�et�q�bUm�(d�<����{s�!M.��@�ɂ���OM�c���/�?��|�[O�̳/�_�5n�w�٧�7�/�m�fj�ˋ+��n������Sct̠}����SF�?B�d"5?���o��d>�Rl����o(s,%�T:��+,����>@<��o���������_��W���_���87����*�r|_5�����Z%��K<���d��ѽܘYS#���{i����z����d�6���
c ��=#,Τ��Np���K�����9�4��D���fX%�Ɩ^ǿ��_c��#�×��7O����`�~��;B2���\#�9�ۮ���!���T��EM|	EzI$\�4����>_7�P����bG�/b����G®m��K�͟d�7��ic��X^�r����z����uU�\m2����Sk��HYz�Mf����������F�� u��4H���iҪ�:�8�M�>�:=��V
M&�&��u����S�
�̥N�mf)Sg��f��ʹ(��M�G�X_Oi+��dUU�(���d5�u�*U�d9GGX^�Q������Z)j�l����.����1_��T��Po���i�w��_����J)��H�ʜ�?����Pnx����;p����S�n�{۽;���ut��3?46�{��<��2*S�v{���F��y�.W�TVf)ٶ��Z��f\v1��v���#d�xq��$*�n�i�Sn��;��ML-#C�����4�n��wh k݁�=f�N���i��Ӄ�,̠���α;�ucd�Z:E�&�b��YR����p�e�nr������Be�"�>�Cʍ2k��PluŚO����enq�����PG����R�cajF��|���4kP��-�`�(`�Tȩ9��T�zUω�>6�UA�L�z�����w�`��(�Hw��'I9��L��W����ْ��R��8�A�܄W�K�C]DW��U�$���t2�藉O�*�La�q��F����-dsiV�W�������Z~J�t�	@*�1�ٓc�q����xŦE΁<���� ^T�c##Zb?]T��z��0���Xel򜰈��Q2npv9�m)Q5��PD����m2!��AfnNi���ng��qج�)�[�6V�����PX�Q�>j�<�3��r�}��xg��1[����[`�3y�*�b�m[�9s�'ϼƶ������S�=���a� F��g~�4'^z����\�|�������n���\�����[��?���[$�^�aI�������_�����ě?�Z-���d`p�T>˅�x���<�:��ض��O����LK�x��6L�d��03�2���6"]a���mu����2�VN�J�
;���&�l���t��1y��ߤ��Ǝ��LN^��A�/̍���q���_�S�����������§~�񱝸�= ����	��B�f��ir��gX�~��'ɶm"�q�X7r��E�VW/.��X"Ž�Od`�+W���W�����������s�,�x죏i��3�?���Wx����'���;8����m���K�={�G�;�ڍ7�&&�e{?�jO��L�ʵ���}�D,���MX��.�����F	��I_��B	Q�b�i����j�@�8��mDe|� �t��뗘�1��f�X,Uh�������c�m�9u��z\���9Fo����R��.��'���Կ���ry�ޖ.��IjM7�?��� ��0+���%$@����C�X�h��25���)g�B*��}�����x��.-C]m�Ģ&�tᶴՊ�dlӢ�}��wؔ~p����B��U�X��&y� 8���n6�BK��]��&u�����y����m��x�
V��l�L�j�+��UNck�}�*��V��L�QӹC��QOK"U.���L8�j���)��kP_ފ��t��J*�\."qJ�5%]�NQ��!Q��u1-Q����W�ڥ��E��k;<{�����߿s��{�g�]1�W�>>~��_����i2�M��RG��*��-���br*15�� 錈QDm�O>W�r��Z$DHʉbr]�ܬSkTh���OL�k�-�b���a~i��.��8d�,g�5�XXӞc6��,YvRU7�����} vN�|�KO)K��W�K��)��~{연�x�~�~�MV���;��gg�"��w�-�LvF�vr���nβ[!�<�h�C����>�,��Ŏ������}T���S�t����N�9e��o�R��u�wl��t/ea��j5�
�{z���#�M<���,�$%�y�</��0L%x@@��_���1Jo��aU`(@F@�� �ܤ�,̛LFr�'P^'�K���Su��S �X�H�UƲ�Y�o�>�²I���x��b/#�,���_���{��fV��rYA��eC��V;R"�q
 �N^���s��Yv�ءc���N�.���0��0�X�^Q�5tq &ދ���{I��X ɱ'b�Zv�����*�^r�<x�>e�ľfU"�,m��,���w���O���	c��9�*[v�#�<O�c��+�SO���7v����,��M{�Z��T?���I�S,,N14������r�b�E�l&��q��8�g��g_���A>7K����	�p�����c�.]�ҹ��IM����@�V� o���<a�M���&�������@����f�?{�je<�,{��a,f�z�H����E�f.cj����6?F�ݩ�DF�����ҩK?��Jb��QҸ�3�����R���{��t�o�T�l����G1��L�k}��Q�\��l���!�����blݠR�dh����Z%���Q����lޱ�Cwը���(���wX�[���ǣ�{�8��9߱�2���������U�����GB�^>y���k��8�sTh/���� �AI��g>Z���
f�G�������� �)t�g�Qj�5<��a7��(�f�`8@��&Kr�ȷ�ή>�<��L<����@���vzzJ$sˬ��<��c��~��O�����e�.?�����9��&�.��(��L�
}C�Ґ/�p+��f�����^^;y���ჷ�K/������"͖	o0���"���Zet��֭.��{o�����OQ�ϳ�M084�����KY��E����Q3�e��,�)�tE�:}����H�
[��V�U����"q�F����"�efv������*��1X}����Q����x���o�����
��i�)>�&�mQo�0�ŀ^Rs�[E�e9]�^s���6Z�m�`~9J"�Q!M,���n�� ��K�X�nǄ�_�L*I6�R0(�PD72���.�F��	�^��[����*S�{�������+Px��?�߼���Kom۳g3��U-͉=G"�R������Z�NLF�6�W�%�M駳�n:��]T**��װ�F�,R,�	���i�6F�C�1լ��1���P�Fӽ:ىW[8�5vn����b3wL����q��}��ߋ�k�����/Ҫ�l42��`����%��<۷����=�}��C��E������r���"5��:���>C!����Pn����ģs��=|�cS��iaќ�&����nq��-��*H�Ɇ�W&5^6`e2)-�
K' �\)a�t<��VY��N@�F�� a���@$}o%aw2I
H�B:��*?�C���>N�L��+`J �x�����'���_��s�N��$oY��������ӧO뤨��Z�%�$67V�+���Lr�z\/��E�F�C������u��s&ۭ-/��/׀�� ����(��P��) PXD	����p(W+P(�Ec[��\�O�H��E�Tya ������1��_'�s��	x\�E՚�s��Yz{��W�	����w���Wy���l!Wʰs|�r���>�Sr�2[wo�я?BUlT�z���y�lv�z孬.�5��z������e��o����gy�O�w� �����\�@�V}��?s���q��C��*-��LY96l�5���Jtu�z���w����D��Gli��~�,����m��Y��q���	ww�Z�I���h�r[�ŧY�^�hv�!d6��]y�}ˣ`qKF%�^�ю�ٶxս���D�FYY/����74εk���|���F������%F��>���%f/6c���|��1/}�>�{�T����������\��J���#���,}�ӓ��Q�e��o�&��%\NC#��sI��$��c��u���'iV-8~�w>G�'��bv�*s�^O���yvn�����
]-�����o+Wn.RjX	���d?�u��"�\��b��(�pH�o�j��̘��P3��n5K�i����&�x�.|�*�_��@蓿�{�ĉ|�{�^��o� �ݣ���2��*���wV�yBA?��*������;�|��7n�&��<�p�����Elf/>oP�;���.Z�K7/c3�ٺ%������KD��ɭ����>��Ӷ����l��K`1�0������V6$�@�v�IC\B=:GJ���eVk����TTDf���.��	���f���U��xl�����#=�+9��:��Aa����N��B�Je�b�-f6��?͚�%̤2��:�t���a�(^��8�~��V5�FE�2��3�T��u�����:�<n�e]z��8�f��PP��nj���}n�M_5>�Q��x��;�����.}{���_~r�װK��ղ��5�D�.N������Z�d�ؙ��V��:%K�]��]YT�W�ģ���D��R8MmZ�
f��7M-~_�=;vv�Ie�\^��2�"[z�
���R�����z5��U1��lҽ�~�+v����j-Ɔ�q��g��\�
���Z*�Ju���*E֖�p�7��7H��a��0�F�Sg�b��2�}��l�1�]G�����F�$��DK�v#�f���~�����m ��q}=��NJ�����1H�Y��zH��e�и�2"`H~��K��L�29��T�h0(�ѿ'�K��� �� �k�L,c��tu \��>��oa�6loN�<�v�ƥ)#���{�G�sQ��2�
Ќ����R� �"\!���zb�-̨���۫�LGfgپ}׮\U�)�/���]�0vrl�O@�<n�]�7Ao���8��Xb��l7���LN���e4Y�I��!���s�F�ĻB��� �
��I|� �TR�*�]����������S��dfy��g�eƷM][����Ȥ�|�|���۱yL��B�.pr�9�zz��/LI4�!�G����]��2���#�#���4a7�(�Ӛ�[7�	D��Ѓ���WN�p�>��mۯ���F�l�lrc}�Ze��/kז����~�.�]����,�n?�FQot>w�l*K:�^G���ƺ�IS$D��74#�sӨ�hTsTk�TM��3��(�d�z~��+O𴘏'87ug���B�b���)~�&Z� =��[�1�=z]D�$�	��d�t��x���s�u{�z<����鬙���߳[f�-��-�i]��w���������\:�_��'@,�j��<A'���W�6��G��/�ׯ���cw����w�tx��e�y�������=ҍ&��y/���g�
Ng�x��r<Ǿ������c#C�Z5��:]~�(W
Ye�%CZҗ$ZW�̎ 8C��Қ��ά��<��`?ֺ���7�2j�i(/�����	��Gx��9y�{\�z!�8r�@Ы lyiA�)Vk�\V���)T$��I����Ǳڭ�|�b����w�����R�ӫ"������gg�,DBvￍ}�ZHP\}�5M���9�^nb��z+�� �ɸ���W���)�`5[����,�QI<
`���aw�l�����?Y�m^\�~V���nr�<mkh��6�B%���SPhm�i�X\6��F�uh��$���U��덖��}^��^�`�c/V�ֵ�p=��`�i�D,�T����KY�\6��s۠���%��ښ
SUE�:K�-�[&�V6�0����}h�?�
��H轗�s�(�~��#/=��5�3�A�F٬n���;�j�|Ro�~6��~54O�Ɩ�1�F4��ܲ�94r��n�(����P�Q��7O�PC_	��>}�x1E[T������Y����G�Y�d��-)�u�19���%�rs��o`��9t�]����
zپ9���3W����a��h���?#��ӷy���Nw���uz#;H'̼ua����=c��s
Xz���N�?x�q-�H�e�`�ڕM�:�1�]��( sy:6$"� �SP#��E�ߓs*�])%	���;*72���y    IDAT7�b:�߬�pI/� Cs6�CA��_��a0](vb�d_�Ϋ� #��We�۫%f�r���=u�NX
���w��2ҏ%�l�ho������lS +l��O�r#�N�&y�0��J�_���`XJ�2^�0L��A2vyo��4ۨWj�)=��F�;'H�z���ݳ_A��ƒ��
wV쭖2�;����I-su:\,�,�]Ю[�������.S7��"��{�E��x�<;&��G��������^���͌�m"�siV��V>3�B[��|����,���vk[������ݬb1I����I6�������,�'���~Dv],x��2���EN��[4j,�����e׾���Ώ`��9��y5��4�3?N�z#C��U�+fK[�J�TҖ��ф��崲�8I������d,3u�)b��K?t����L�?��x���R������B�H��P{�f[��L������jE"�J4UV��z����Ko1y�5�#a�����
���/��?0;��~/����1<�o0�g9u��rA�]_���pW���y̶�����$(
�XF+%���Oaw�{/s��kH�2�v��Q��,�������2�������E�mS�����L�h5��mF��"�z���AowH��d�g����"2�ϕ�X����\M��K�Qa��������9|��B����O���V����g𹌤Sy�>|�}��&�D�^��S�Ӭ%r��}4-6�Y�{����G>��k���7�F)���Op���������gv~A�1����\ۍ�	�٦	)��ا���L]x��+ߡ;(L�E�;R]�Pf�z�ES̠[�Mq�h��[@���Kěڴ�YVM2S�;2J��,ڄ\hMj�/�pe5C�,��!*Y�.e����
�DĎ�^;}��V���HY��Cc$��4�^��>��s���0�f�X�5�(P,�`Ȍ�h�e6S6YϥhK��Ԧ\+����R3�]o/f�`*U(#V����;�]�cv�2�0Z��8���Ờ_|�|��{�g�]�����F���޿��Wn5�
j�i2�Y]6e�lv�^���$;d��<m��q�f ��a�[;��NY�>kU]U��Y��!f4�d8�C��E��(����ڿW�1Q!b��k|�b&���m�f�2&���KTW��ע�Gv1����W/r��=x�C��b��TF�?d���r���91��m�"w˶���|O�E�XR%^�R#en���T�g�W߼IO��=���&�9��>�A�;r'_���� L \1-+]���PH��L������HDmغ�' .�N��ۧ��RJ�IV�b#�x21v,d<��!�^'A�:o ?6�x"�! M@�����3IuZF-�������WD@�Ύ���%~�R.���"����,Ǐ���G���E�m�D����w&�%,�!�z2&�˩���s���w�u���ޔgg���Vͻ%*�\ֱ��^J��c���A���������G���6�JI��ض���{ֵۨ$$���������w)���r#�Uz��U-�����<s�S�rBD5Ul��p���v�؍�dx�|�䫸6|>3��,>/]f|N#I�17i[��(�?F�X�n�j/�xمN2�8�VK?#aZ|>)SՈ�ʬ��{�p�����,��������lPy�0��k����	vK�������e���(�7W�y��&ƨ֫�t�5U {�aN�x�)��ҤV�7�Y߫�4�oQ6x��%ξv�����Ls��].���|S�^��Ne�yL�$���S+�Aҥ��m&2�k�]�`lzqY�ڪ"��r�Ǎ�j��P��Itq���~����#��u�{�G�O���j������g�1��n.]=�?z�b9GW�x݉�ܲF����KD�t"Moo�2;�J��>�a�)�֙���|�Ng���[�Y�E���`�����	�YX�2f���*�TJ":���L�vE��zE�Ka��!�R�J����O�.�A���݊�ndu~
S�L���FYJ����ا�<�MT�f���/1;{���F���~�F�E�X�PL���0�̬�p����'~�CG?@��f=���W�gea����J���YDޜ��ih�y�(k�4��)n;t7Ǐg���+>w�%�?�?$�H�M5����e��jǊ�`W+ sӤ��l�k�����&�ee�EL%�OC6��x��p���;�,���&G�R����b����E��ҖcWEvm�>G]�
���������1��F�������8[�o'�ɓˤ���c�@C�5,&��{SZo�iH��H<����l5RoW�;-+%�r�f�;��RZ7I�R����l�m�Rm:������/~�=�ɻ�D�m��@�0�?�֟<yp_ߞdv�cX�k
�2�?�����ZǼ��W=��ԓ�z��ʥX�N5z��x,�Z]�(;Qz�ʒ��WձX�����Q���ϭ&XI�W��(`i���y�i�]�V�Ѯ��%����bo�_�b��ʅ�5��دQi�������P��ٓ���qTRx�&��;v�"�q����6�1�N �e1^�X�`�sQ�%��F��8,L�����w�K<����x�-�6_I��ݯ��b�-,�4"�A5+��0�TK��O^"W�]���f���Qm�exxTY0�,�	�Q�0nR�%�0kނ��5��	�IF'U�Q�I�펇�0��S��HM��uۥ�Q�	�M_.(��S�Lz����������^W�N ��D�	`�PK���C��#�dW���VhR�Cj�´��I9Y���N�)c�+�X�,�ZF�hֱ�����fK�;=oǢ�A���	�nJKC�|&Ǧ�q䘥�����g�-dɗ��@U�¨*��DX^��C|��w����({*�N��r�4��ĒI��:���+Wo0=u�ˌ���aK�x�x�F|v�|���籇��~��n.�y�jr�ŀ�]'�S)��#t�q)7�L��H��[!���x��WYY������N��c4Zu�B4꫼��?c5����B��>���}�L_����]�L\?�t�{�y������묬��{)�2_H�����[0�-�:�s�np��[�g���y���������n���V�?A����j��W�;�I�`�b��YO5q��؍��Y�c4H_a�l� 63�.s�7�'���'~±{>�G�5*-+�N=��7�h��Z�N.Q�Qt]I�?<������z[?�f��z<N��K�Y�l��J�+������(r*r�����B�+@=_�`�r׃���%����|���xD0����I-7���'�5S�)��\SŢ����+Y�M,ƍ�L
��I�։���YY�qtK�����J	���Ý�|S�Kj-N0l�v�so<���yR���<斓d<�m�О����bx�n���&W5�Lg����-27u��NaʮbmԘ�[���Ȧ!m�1�Z��>v<��=�-��ᳱJ��sdN�d5��m2���djS��5_���x��WW��;s�<o2���A���e
0b�Zij�!S�u���P��8�.7͖D,�}
���b��[\
�52�aK$���"d�e���i5!HoO7���X:���X��t���hsR2���"
fa2[�VJ��8԰�:�Qz�u�h���$\��6����,�6�p���[�|��߃6w{�(\�zf�Փ_~�^^9P�Uٌ��Y7��T�
���vIA�0,�]�ۈ.K�oC�:�,#_�T|�M}a-u� Y M����O�L�GI��r*C�	�Ŗ�~�QF{�l�]��/����|���+9�l#�A��k� �__aﮣ��ޏ�tbqy��sjlz��k�ş�����V�##�t9xz|vB�:NS�R#O��Iw��S��5B,�

l�����ϣ��Ͷ�����-!�z��j4N(�E����rj����2ã#* Y�Fٿ�.\������X��ϯ��7�o2�u���b��x4)8��.�������L�L0	�ڈ��%}�=�*R1����S��}l�p�x�u�$Q)w�B
Ƥ�+vB��!�����?� Onrʸ��
�JiX@��-˸��~-o��I��<d��c����"�
�)Y������.y^`�VR�9�0�ּ��j{u5��9�vGp#����pO'f%�c����I:�Vt�.�yI��%��ЙZ��{�~�����o}n��߾��޼u+?|�ǔ�5\��ZP�m�~�'�|��!�����ܶ������M�a�inb�F�Рi�a��_%���O����1{�]>\�6~�K����ЬP-�1��X]�T�=�o���Z��~�{�q�CLNF���9�i,`2�X]<E6�@0Ћ/8̃������+��������8�R��;Bݎ��"��B0hE�f$��dvP����%�p��+
�x�&n\�H�����"V�.?��#\��B+y
���B,ϕbs�TmPiWi�-�+,F��7�s�05�<n�Z��IFƅ������R��;�q���o�6��_8���Nzm���ksY-	�(��uP2���tSn:>��(#}��d^���~V�VTH�h�����6(ƶ���A���c�&|�!>�����'*y^9�S��I�b��9�2�$Q#� F�ƫuj��.��;.��f�&\���;D�g��W���!�<�`��Ġ�;Fp��Agh�X���ə�m�qR��My�|�i��)�a֖�x\m�����!B[w��]�����"Q
�9cQ�Ĺt�F�L/����̟�ʛ7�m�^l�A��y"��95�2�͟������Qm7���(�����[	F@'���~G��!ai�yۨ�cO�i_Cii���|���	h�9�

U䗭���J���N���/��������^��)O����S�B�B�`HDP�78�yu�����Ɉ��PK)#r��y�,�e�4[�q���6�V�.;�Z	�]�-uD�	��U�5n�{��$#�ܨh_a�kf���{۟�gI�n�{۽;�«W�q�{Ϭ�_�q��}8\=\:?˕+�:��vh/�
�p�nan�|.��Ф%=�UY$������7��c��,9�a�n��D�Y_���v+Ș��#;�m��E�>Q&�/�R�ٷ�	u�ʱE�`��� �b����*a��a���)���Z��,������2U0Z�DF����Am~1(ͬ�2i��H��z��K4)x��d��TZ���Ƒ�����wp�ჼ���H�b<��g��0�)2�i�b���:}��i�c񞊮���x"���Mg�I�T�VQ��F[�k,
�6�焵�^=YM� #��)�&`K�P%%ka�TI�߯`\���\.v2~�	8ܰ��'`J@aǧP&\I�)(�}�~k1ݧl'���R���. N�[���0o�2���'���ݽ
be,R�հ >)�ʘe�}��e�����Sz	e���@�!`P��r�J���]�C&�U��ǔ���~K�Cɵj'I&�ݣ�v��M
�žhqa���.���4KV������X��7T�}��1�~�Y����.IoQWW7]�O��Ǹ|~|�=ܼr�|�&G�y؇�T�o3⳶E&���f���?�,6�M����Sw;i�3��.
T��(�A���J��j�7w32q�����}���A�3~�0�&X-��yΞ~�Xt�m�n���9x�C
���os�0�l߶��?�0�\���8=9���R]u�A������kW�p����}6b���\E����v�ta�q�Wޢ�����:צ���J�(*"1Ah�9�k/���1D�b�������l)�?bc��eF��n=�A�}�1-��6��(���KS��1Lu�V6���lٻ�T����e0R�%���]lk/p�� WI��y��L���l��Рz�Z.�6;��dd|/��G-D��klJٸɹ7_�ƕ�$�+8�&2��^s�F[{�m������Q��&ʹ�Jc�AM��$j���*�@���p7.sCc�zt�og��%�}����}�6GX\��2=}a�]8O8ԋ�!��d}�&G�ަ���k7���{� �������t�yr�A�I ��i�"%*��V�-[��v]�l��V�u�׷��{����,/%J��HJ$�b3�D 3 f�g��s��޷1�����]55�3ݧ�9s��=��>��R.Wu���V�`%�F�,�~�+�,-�P�A��8��]�~�e�Vs�N`�Z)����'�F��B��$S�i3��.sX�U��I[�rn���4��:/���W��|S�~��m4�U ���²iU�ʘ�4d��qD7q��;���C����U���{�[�S��H{#C�0��.�f��i�s4�W�x�b��S�Q4��1X*Ҩ�
�W.v�u�d�?�J6E�ja=_Ԏs�S�]J���#����*m���+>�l�[�JM�ٰ��V��s�64-q�l��;~��|���:�{�g�}1�33��O�����խ��f,F\-&\N?3W/���%�_`l���x�p؏�%Ba��2X]^�)��p���Oji���J6���m���Ŝ�ܵv]�����S���Ud�k�k��v/.^fznM�Ⲋ2�&�ܵ�b2K��Ҋ�s�GX��x��BԾ�H�ȥXKNR��cZJj=q��{���>M���>�Y^$�3�:-�2muG7�L7���[l���[N~��OU/����mer����&�?p��|�{�8�}�C$�*��Z�h�[��/ �TT�/ Hk�#,��׉g�wQ(����ۥ J����k�ϵ�FO�*��,ڛ��Pe���Q��*��	x�f`���w���	�'�f��`)Bh�����D,,��`{�]�\��Lf���ݽG�)ǐ/4�[����q��CW�E�O6��j��l*8��%YE�Sz ��;��6z���ZX;��싔wŢF4�RV�G��=uN��Ĩ�@)H���޽Ȟ�Q,�YK��r�eL�f���er�Ieze���7���m��K��}��|�W�~�o����\�:�y޻w���ko)��e�6��e�$�q��A�u#�Z�����xI���F���R�ۨ,�d}�8O�%���,H���a��j�� Yv������GX�:y���[�F�ak�I��	�<KWy��o�K�06���|�+��#[�������%��b��D��������da��r+��W�*4�]�>�;}�r�4~�>�˓�O��H̅��b��hŇy��鳯�u6YLWy��E� m�F�RQ֨Xlb�y�i�����.�N��+j��3�E���Ũk��c�=ŭ�}�>�E�0/�&1}��ׂ˴Ь֨��Ʃ��D6M�o��%�j�FXK,�q�iV��n,��L�`(����R�j���ؒ���-�ٷu��������^�Sʥp9��:u���I�=s�R6���'N���{g�rEw�ArS)X\���[���#�+$�)�����s�����ai��$�pګ�?�#��*��͓�r���M,�fu�*݃q.�ΐ�K耗��G�T��/���u_�a7,��#�qY�Jբ ]�`w"Z�����盔%�����h2wc����V'�\	�݂#�V-46;�z������V�8%���m�-�Ҹ$V`��I���qŴ�<["���n3�TKz�ʽ���R�����{��4���Fԥ���z�F�FW�&7��*��4G��
5Cu�MC|.�6��|6�&�PXB����)vW>�.ڥ�D�J�)L��ZUZ��'�~���4kŴømT����P*�t�����o���f3�BVZf�Fۊ�����������f���)�\\?��3�@�ŋ?9�ҷ�����f��ћ9{f�w�^f˶ڔ(VV�x�$֖銅T,�J.qg����ed���Y�l�N��aye�f#C�ݦm��)��z���ҝ�g1�&׬����0�QL��;YXMQ�H��T�a7[�xi�ӿ#W��q������ȉ��A1S���.���<s��4��]q��?��+��_$��6Aw
�Y´ٙ�_�����*'OU�_wiy�Ep�=    IDAT��Y�<�����q?;F4{��{?��w�����9u�.�_W���"���t) *W;^UWff����h�t�s8t5-:0�h�U�0sL��e��C�k&�Q�! M}�Qe�X	��FYY�������P6N�m��E@�����iF>�o���n[ �lO�/�V���d���N�^]���E��-���1�<��aL�6�9�'��:��+��<m��Lj��ի�)�K��[)�#�&���j�9�P�X�.������������2��$�(WK�%V�Iu�6�)�c.*�����-���{x��S<����۽�b��ϟ|�`XJnYe��GF)�����.�������y69�1�`lȭ�Í�:!��dԩ����ġ/����OH��a�`�J8|��4�݂�h�l7�(�jS5b�#������u��mc�Um����4h4�y���)R�����}����4�N�Ǿ���'W@���q��X����gĬڡI:�R�R�vm�Ҡ�/ν��K���/�oع�Z�`|�^�=={�i�۳��u�/d9{y�/��>i�r���5v?cC�	��8,�,�R�)��Q����������K>|�op��'Ul��?`�����6����� ng�F�����JN�:I8&��M=�X�t6����em
��e*Ŋ�ǘ��Jb��r�R1Mnm�#�������ڶiD����o9}��VI��&�]�?{���͔�b��'^_����6	�.�\�|�hW�\&�EʎV'�Ƿ���:��	�.�r��K����N.���x	ZK|vҙ�j���AV��0�C�b�߷�奫D�M��i�J��>r������\%�(ɢ�ZI�T�eW&�T���C��F%E��Q�S�/���g��]��n�h5M�-a����Ь�q4e�%1�i����9���t����qW'=���]YT�t2�k

�:���x�آ�h��	��#hU���.�jx�������XP�gi��p���\U�����ʘ"i-���f���vǛ�ݨwJȆ�l&׉�Y]�h��,:��*V��P�W^J�:.�Ĉ�4� F��P�T��:��� ��۱� ����p��?�w�+�����w�(�·_�����h�����S�8q�j �������H�V�����b���l�4������Y�~�j��������X�z�t�
}Q�ں�[m���kHvy�
�c1B^;��t��XVM�r�N��U�i��~3F��:|�;��ĹY��Ь4������)��f��{o�#���A/W�|���I܎ꍔ�V�Ħ-R��9�˫d�]�V�l�w;�P7�� ����w������_�W������7af���m��� #��V������e��������;+�j���b�,eUn�6��RBFPJ'�V�C��>T�9�����O�
;���uL��CXA1���I)I�W�@a	5�����RI���N � =ٞ� �'ٞD�	�W&���� 9\���g���Z�J)��,`Q����NQͥK�ZD9j�c��`�8=y_W� r.�Y�A@����UfNlFĎF�4E�*�t�K��D�{�]�ϛo������ܱ]��#��&�`���a���G)���I)��ؖM�����F�����c�P\b�X��X���Ȑ�Xԅ���ժ��ƃ��\���w�[�^VN���KG	�+�
*�$a�6w���I�-�g��%�5���Mw�-�y��������
t�O>E����k�3?w�;��Я���Xl$/����+����eJ庚�K���¼ZҬ./h�H!+��G�,~wN\��� ��=�$4y�8Akk����tm�G����#��SX�z6��؅�\�[�Nf�4�n�P��6Nvn�	��M� F�^�����K�1\^%�����Kжs�_d��0�a���3w�E��߉�>H�����{tb��r�L�W�-�N�(�x7�B�S:>�z�}�.VVq���$���T����㹧�᪒�,s��q��*���9>p�G�w@��|�Q����ۗ&'cdxWf41ƮF����ۢ0W���me׶	B�&kҴ�����}�KN��{���i�Κ��Z�Z�:�Z���t8��j��|��f�k��h�%���\�TX�]k�ƨ
���gw�X\Z���NĜ88�h٩Ѳ�&�Z��r�ղL��ӆ�֢e�bk�x�Z��)z���~��E�B�~�`:ȗM�WR,'����VI6��#��в��V���7�R�)������m'>o�`$�Z:��U�� �\��n�4q4�8�m-�>�u!�@��*sj:��S�sٶ�bWJ��Ī�Ţilaeq5�ե6���z�zz��\!F�'�J3Q0�U	�ï�(S��P-�)�D+�^m��U�j�ִب���h�����??|���:�{�g�}�B���|��/�Ξ��{�>re�.�wq�����N�!��=���߃)^S��|I�7���zp�xY�1�D�x������Y���"�)r�"�X�������wE)U3tu;�����j�)�Ձ�������V�Z��U]�mwbV��Dv��o��g/�����L�������웜x���.�{�|������?�����+�f�R�И���	�-���㸣;�y����	Gz�8y����{�{ϝL�s��o���x?���H![��g��գ�(��ǻ	�
�d`@$���rk���L��x|�N�E��웰<��2m4�lX�(���b`��q� Iy�zӼf��a'�E����i+ݾ��
��;W<�C�/��ȓ�fL���,��j��$E�-�I��g��>x=��=ٞv5[ee���I�� @�R��)�S&#c�͍2��F�Í��`ʶ�'�CQΧץ%�l&�̣���fZ�7Q^/�����U-�z<n-��A��Wx��0�y3���>{���~����������Q�>?�G>�1.\�����1>���.��W��[t`ej�i&F����
���J�I6��c�������t�z�2�4(�8=~��	ݮS/7h>W+/;n�(�J����А���,=�qb]Q�'y�'H�/082���ؼ#x�v?�ٷx���=����Y�^j���<?�8��!���g
���p����W����N������o�va��3/�.M�q587=M|t�b�����s�-���8v�"���Hf���~�V7��BQU1�7��y*��iΝy]����ax�s$3U�߿���qv	�����308���)~��o�I��E���%�⒔b�&�b�X<Lbi�с1*�6v��?��?��;3���S?���M<dr���y<��g�uӽ�Bc���;�IV�f�1B���mۤ��co����@��ڧT*��!�������^=�����%f��9�vY��{�^J�4����*}���O�Cc}67V1�2��Qtw�ȁj���ō��ZI�j6h6�XM�9�;b����R��u��.i�*�Kzݵ��n�q�T.`sش,[+w�+�]R����&����e�h;(�Lj��"�1
�A�j��N�����dK�2��1.]��>�]� �Z��h�j�H�Q�B�)ZBiL��*�#y�u2L;�)�{-j��R�m�ak�VY�>gS��m�l��,�e�TPOHK��!�&�q�c��ޯB�\�EtB�|!�SY
�6V��t����f˶]x=�Ʒ05u���1�p�F�$�W�eRˬ�^��#���wRy������l��4��v$vۗw����~���]?��|�ѭ��_���0�o���'v��ݼ�����X�b1��"ʷH�I�B��#�X�%�f�n���Ao��$ ��8-��j������6�s�I������v\6Y�Y�ԛJ��mN�ۦ�z݆�*^�bZ�aqo&��!�f/'N��7r�&�ʩ.I��W�N��K?#�Z䆛n��~�w�f��~Wm�R�,��;D&W���s�j�׎%Y-X(�q���#,����,�}��z�l�8���m⏿����-���o��G����������5�z@ʗv�S���lM�P�&�������2�J\ �<���&L��$a=DɄ#�I�@2�lص� /����4t�e_��KJ)׶����~���!?K7q��
(E���T'(�/�"J��ZN$Vٽc'��=��ny�믽� R�K|n���vX?y��ⲂC�Lَ�E���S�;�w�6[(�k6i�1��	�OȒ�ZM\�����
�E�&���u{r��d�|!K:��d	)7���ĦM[��37�c���ƞ�K3����CC�����d=�f��=\��兣/3�?B�.��i��&�>b�~#�ͻe!4���bx0�H<Dn=�����C��h��.>���+ļ5l�*պ�i��/����a��^o �+B��$��˯�R����/�6�[���v�s��������������,�o� ���?��Jj�`��ۯ?ΓO��rJ�*�J�i!��`���ԫm���z�X�vK|��c�H<Э�_| ���}гVR`T�:���%�nXJ�10��t��R���|�������l�m{��;L��PP��X��jbw�XK$u�<y�e&/�B�碫{����y��%^y�(�\�H��g�-Ƨ?�%���jT��o2;}�J)�g?�/��*KK)�(�v�Q����\��Bb��@�я�
��̃�����c�H�Y��X���-_��M7`ur��y-�޸?�˜;��F�i��Ң�wǥ�#�{¶
���G�H���I���G��b���ꕳ�t�h�`�jaumW=���0�j���-�aԫ�~��eU&�\nvr���gP�I�Z�o9Z�ng�2l��a�N�S/j��b�f����T�ee��N����{��H�h{��yr��g[[�o�mUq��T�HP�Z��q-��U�{�ٲ�)KL�U5��H�-Ъ�K%1-u<N�{�P�b6@!�

e<FO:��59�؝��2>������U6�G�fW�ċ�hc��0l�Z5�D$r�Lj#>T�K�&���ua���1�zG��"��ӱ�P�؉IEDt�Rebp��Օi�볬�L24#�6����q_�Z�Z��/p�om��?r�)����x_���ѯoK^��K!��X� !�~�E�va	���� ��ua�
�|J.ҙ��E�u���}j��5\�C<��c�������m0�u���3$"0�]�m[F۩�S8lVZ��,�ݨ�K��ϩ���j3M&�����vNн��n��:�aa�[Y�B���m!�����i�UP|��ڻ���ӧ����1)T*$��^�	�M<��,��Pjy�d�������G�C���`_�c�Fh5�ڭ�W��_�V��^�#�0}y���~u�����R��t��>�<� .F��:6-�.�6�s°���4��0��dR� JeW-�\K�}��P(��L(R�M$W;>�m���
�� :�b�#����7(C8�e�2�/��B�Y�4����[h)���0�,3��)
0S͝˥���"i��F"�/l�FiZ�Q�6|��;M1���z���j�F�8,m�v�aw#�#)�[���pIrٵw{�����C��]:Y�7g�TP�ϑ#G8��)�� ���1=s��v��x��7�1Ƀ���k�o$���3�G��L6�{���b6���N.���0	Ķ��_��0{�0k3��汶�4�6*m�t�E�feyiIb�o�p����W�2��nn���hZD"A�e�~C�b{��`!�"-��{?�km�dk�L:q�\1����j�~��	V�.S�%�;����tH�*�QoH�z�m�lr�>���h�
�
4�Gq��d�K,/\��P+牉=�J��"��l��6�8}�<k�w|�K��;�U6��{�޲3�y�Ο���`m�$���X�M�vjY��ɋ8��ܸ�N��
��'��'����i����&41���7���O=��[�l���.���'�_��_�N����������	K�^x�Y*�U�d1V�%�Qw{ؼ���8?��a�m�n����%^{�87�Uū�)_,J3�M&�&)�2:��R����y
�%j�EvuGY�z�ư֚6�x�$�r?�}p�m;F83�6v�o��g��"�_�a܊�v�+��f�vܶ(͚A�^�ʏ�~����s��((��h{��[eh������䫋��,JC�.�F�c�Xkam��5���J�Iˬ�^�-z���;�YD�U�ї8���E�&S(���Cbu�tr��x�Z)�ݔ.�S(�P�m��i�-�X05�5mJ�ŧi:�k�!*��z֭5L��aS�_�m��8�:�XȪ�\����3e�i��!U����..N�SiY1�,� ��[q���zs���M�ff��t��2g9���15�.������v���?`�2DBٜ�U^5��d�cu���=7�_��)|������(<{�������<X1<���'�;@b�����Ew"�:O��YZ�Ҵ���2��O�|;=�}����hYZ�H93MĖ#0��afq��dN�zk�<{�O`VS،Nt��BxNjb�b���M.+]l�2%	�F��O�5Ax�C��)r����}�}X���02:�Zb���=����ޠt#&��p�����&��KxM�X�d�جN'�� �+��W�{G�K�4�]��-i����4�j����T�;�0(4�y����w�P���7ayqE���y".��'�&��jgZ:�Ձ[@�4بEL�_��0jr�� ���W�PJ���t�b�p�5_����eR�$oyl����i��D�h:HY?C�� 1������^����n�ʤ���m�g�R��D�NF�`�iE��چ89�n@'��fg4T�(ۖ�j�"@�\��BDH��0�iS��]s$m��'�����!��d�J�h���e��;рim6V�@�H�ݻ�34:̶�[t�^�_aq~A�[�_:��}�+�8�v-A_�<͝w�C�P��Çcdl��g/�y1l-���,s`k?Fy�e���	J�i�YRB���!����x|Q��z��/��k�F�ަ�0�4L�>7��n�|U�i[�l�p��8uj
�3Nt�Zf\���%6����:�2���[�T����0�"=a���}nW����4��^{���.�M�0�:6��L����Z�s��	|'T쌏3�9���1	(���N-M��,�s���H��a�q���o���b���:�|�+L���]��;n��䥣���u��C���v25�&k+Ǩ�Vĩ�X<B�\���y�zo&Ҍj�ʞ�[�������)��Wq;=|�_enf��~�G��_�'��γ�X����W9z�(���Q�'_ðZ�t���������k�̝��7�2�Xd�M���_<�2]�a.]Y�Ѳi�Ķ�{�)lr��J1E$�Y�vh�-��q���^8�h�E�.���8+8��ui��3顒J�Dc>��e��"T�)\һ�w��.�j{��)�݊ѦVɫ'�m�lTp���4"���ۖ����8��b��n��'��zS%-AxMTmH2�m�;.o���梡�--��Q7,Nl�C;���S�g�
�L'=��2YR�-9;��F��}.��_@a��D�G��X������Ѣ��;VR�Ue��6�Q��k6*8%J�"en�fQKVr'�I,�L$qI�G�c�ԅI��v�;�\"�Ď}�p��v����O����apxH5�҈�z���LC��ba���>�L:s���$�V����p�6��\`n������:(����x_���7޺r�#�Vj�T���w���V�e�2^��e8��-%g)����3\8{[��]7�h��t�v�Y�-,�:%K���w��U�OPkUH�ku5U��"�0qٛ�[%��j��:	bf�.v&���՚%,�a��Ph����	�_H�^���g>�'�Ymb�v�^����/~�0qw�̓z�>-��D/�Nw$��cCq���H��T�Ҫ�g^�筤[l�ݎ�4��cnvN��t#�������;h�Ϭ�O|�[ZL�kI�����<9V�6�������    IDAT��UM< &��a�T���`��=W��JlVarN6<ա�:��No'�M X8�Ɗb>��~"�@)�MxRM,8��T*5]#��W�'�M����m ź��^��²��#�HCA���{�:;��t%�{��~baE�$ O�)�%��(��սҶ:���e4���*�@��$�|�S�Bo?�띲�4��ԼgXA����𠲂��å%��Q�w��#�j�!%'��<��TZ�x�?~�ՕDǐ;���s�v�9x�-�����%5tvJ���-�r�3�/�D�{�(��4��<w�t�l�i43�F��A&������Ϫ��ҩ�SJ�%�(cix�������sĺX طk'�P������P�^�6�m�����:����^�ֺL��D0h'���]?��mae�w�CvuA�""���D�ҍ�s�y�G��zC��F��ݴ�X�d�H�G�'�H��{*���a1�6x�\Y�i�p���%��x�3��7jܼ�6.��L��{ׇ�Y�<{�y<.��s;��G��,:p�-���?C�x�,�rI�N�8α�.02q��K���`��eҹ5�x�	-��!��w�_>�</�|���w_��xDsz����{�҅y�q��O�-c������h���<��c�Ě>Ϧ>aO��z��櫧Y^XԜ�ŕ,3I��9@(�\Ȱ�8MM��a�y�(Ȱؽ�m�ܴ17}��c��n#�3u�%FF�8\�v�Z�B!��w1/�ױ5Z�".�� �!ZU����aIU�w-NO��0tv�S��$`3D�XS�{�U���z]kεD�������Vg)^�b�΁*��MK�Y�-��-��ځ��4[u�X�=٨��|w��,�$5T���v�JJ���ܧ�s��l�:�d�8�d,����C�æX�4�(:>��|Vm��u2�I����2nHE@�G�ŭVg��ڶ����;S�R�`8��<s����ঝ4	��DYXYU�����7�o����ofzV��UR�s<��O駻+���Ev���̓/Na1r+�lTZ��=z�]���u�������}��7�>�mq晧��P+�}�i7�$��m�Z,���,�YX^�̅㸻�����D��ϖ�>2�E,f��O�Bw(D4$�H��6��Mr�n$�\!_+�i�4Gr� ��2-�zÊo�;���.k#@��m1����S̺�K�m�o�"��Y������մ�l�J�f�X-�M�r��ψ�	n����`�ťy�|�<�`�ǩ�c��T�E���%�n�8�����:��)eRD�^��=��b��[8��	���S�^���.�7�ٮbdm<� �vlW�h�q8��	u� %^�::iwP",���e�Z*(W���N��oe �k�AgP�AL"�s��n���W�ggf4�Lb�4�����v�)}2�ZmZ��/�ϱ��ue{�p�b���n%���H��Y�P�`7�z|e"%_U�b�8��N�U���d���d����=.m���_���9���7���SJ�b��#�(y.�46Hi���_{)�h�u ���;���z�p4��q��D�K��A=F�n;���I��jM5���,�ؗ��(8�}6qdd���9�~����D����ϕ�i$�/�.�hU�P��;�`�̰{K���Z �mUVV��7v;�|Q��^x���i�����P.�z}��vVŴ=>�@]Ϊ��/އ���8]8x��i�=Qj"'h�����|��;���&�2�D�� �/�,.�0Z�--02�K>+V#V=��LZ��� 9�n*�v��Z�`5�%��X@ɏ��9	x�/�218�˴S�䴔f�X��b�<��J����.2ټVz�C���[��1V3�7_*�V�+�)љ&�z�@��ɷ��T�A,j�:��~'�+�}z�R��-����j���>�)W�y��3<��3,�-b`��������2Rw�}_����կ~��;�y��21��˓S|�cf|�?z���cA,�2aW�`s	G+��p/����;�[+�o>�Gx�|����\��gP���Ks���0�5��H����jۤ޶3}�}�6�7u
Xy��/ؾ%��j�et�@���*��R�Bv�����&�-�
��@�9i�|M�g�D�)�n�Ӫ7�4;��ح���2���I����R@���V���uF�`o��e�h�DGʸ"�yo�GU��t'ˈ%�æ��Ja�(��jU���0�"����,Jd�+�X'�3�֮Ep
�Ski�;u<쌍m�ѕ�UW (�$�C�����c�%^�ͺ|F����ÆtS�.�\]c)�g`|3�����>ff�h�V�z�|��#0��Z^5��^[���+D}6����ƕ���Cw��p��F0"`~�r5E��q�0=��n��R������SF���~��g�}���}c��KG����e���OO���Y�*P�����C6�eey���8ݣ^:z�+R~��-,�]f~y���nFz�(�K,d�t�SϤ�Q!s����j�8��p[�+U�"��:xI)WC��H�������;�b#���l����ɋ�.\����!��<�Mpun�Jq�ve��vn祗_�e�=���$�F���>b� +�"��q�'s~�
��;X�ɱ�qV\+3�������W�2=������v	�����t�"۷o����c��qp|�0�D�B��:��Մ�_4�WπZE�}[/Y��j�T�4�h�ijtC'(���,�0]�|As�=^�� UJ��b�,�K�X�jS�_�VU�F��*L�J�G�ô�;����ue
��ްR���@�.ҕ(���<ZV�U��`_�4��-l��N���LT�hz��<�q�����]Y���r_�Z���9����.�L��(@U���m�5:^��˫j�-Z.���Ie?Ν;�������h�k�j�u&�z��n�k_��^�d��e
����E I	�t�`8@�pӳg������-�<��=q�6d
��a��}�P���SO��z�����]R�ܐ��zo��ׯ׀S��+I��.�aN�]$]�r�?�����:5��5]d�y����JbY�������)�h�:��D�4�Yn��K9n���W�߲�M�TՄ]1x�ڦ�\.�vnk�hȭ�,�p��d�X�X��-k�t����f�M���՜-B|x�+yܶ ����Y��E<}~����<-C�h+��D�XZ6^8��#Ll���\�ށq��AY�������q��)������?��/�c�6��z�'�ʗ��`��˗�v��я�����9q����[&��ޛY�=An�$��N2��w�>z����s���/��f�%��y�^��#";Ьo�2vV)_Vua���K:��۶�ie�i5���bs 6D!5���똭U��*v��� ׺t�
5&��(T�$z�k��T-dq&��M��$%���* I����M���|:kP��(�Q���4��V�0�'�Sr�;�P�	�� �el�hVp'~}�6��;�5�'����O����;��{y��N��kU
�.�P��y��Qy�\�)y�m�Փ�r�w�O����_���ȔC�-zͼ�o� Ū��34�~ܡ^�ږ�����Y�I���[���F8���n��Bn�nYT�+L]8Źw��lI�����K��U�IZ������~���͵��;�A�	]�{g�}���KO��������V܁[��8��	F���uSJ��p�-�<ҴP��;o3}�-ʫS�������hT	E��4�����C%~U�F�@�$�2�Ӯq���dZ���s)mL�ZmՠH�X�kL\8�"ۈ���!�ͭr���j)m��!���&X4yba�K�	;�P_疛odfz�lт��'�I����J���ǩd-E?�gJQ���j�F�I��e����[�m�F����,.���Z��7��R��+�.29�.�6�i<���7o�B,�f� �r�@8@����*(vF&���M��R�)��ܢ��(&�� .a$.�X(�K�W<����&
y�Lw��C�@����E�;ҩ,C��k�\^��hj��#�`�D��Z���lK�.�ϥBEu}�o*"����D�DR�=a�JU��iBD1�S1��W�mX��:L_�v��='%��\6��eҒ�EνL(�9��N*�;���%�e���Q�6b�4#Y��E�Ʈ�XH���A�'6)����/25u���MʌJ����T���gs2{�2��(�s����x買ػ�����vu�hX&p�2�us��ݟ&�a����Z+��X�1%�b����z��4�\�X|3��ϛ�Or�75U��2:>�O~�8��ED���8dh���o?H4���KO��v�����62�èW;%5�j",��FÒN��`�)�l����@���'5�brݠ�,���T����?��j�|Q*���O"[�����x���U��׿�K�sTKb�_�4��MÎ��TK�-�c؋�xX[.�{_��ky�֣D�"�o�IW|S���~��s��c>r������;_�m��y���;9x�!N�x�����"+�s�o��;?x�/��o�L��|y���07��c��[��N�������3��d��k�?��7�b�@.�QN;Q��,����L�oY8�e���lo���q0M+o���=�yȗ���:�ڕy��N��fz��2�����K�1hĔ��
�4G?W|e�%��-Yp�*�*��kRR�t��,¤�+6-

Lm *UR��a�dѯV�טCe��B����R�mɾ�=$cZS"���Z��FԦ��{ʥ����u͉A@�>zc�,�\iV�ߋ�R᪵��*�pz�^����hY�S:�EcX�is\s)�M���jJ* -�G���I�����n_�	>��C 6A��&荪\F�/!5H���8�^�f�������e��tz��D(,vBil�v���#�wǗǷ�}�z��:�{�g�}��7�|x��ŧ��WW���ch�fƷ?��IZq;\�^�BW��G��-n:��X����!N��$W����Mͯ�%F$P-W2�UA��K,�J|W$�Q�{[J-I\S� �a�d%�ÅŴ`w[([��.��N"7|��z���eq~���� �Ҭ�R>���)[�,-01��v(�o�^.��D0�!s��tZi�d"K�����>w�E�8s+�b���a��i"�n���ω�o��r���ޯ)*K�	��&����S��(o����$�=�u���T(G	x�Z�rEC�zKS�NdҐaY��@�R�+a�d�-f�j��vn�O�D$���DXy��k� �NV�:�V+��HiV�Z]��Ѩ.a��l�9�v;���~�0��#2�oD��dT(�p�}:(oD�IS�he ��UK�$���\,��HR�I�^��b�X
�	`�Ք�NXGy�a������X��S�s8�s7=;�:$aMW��T�.�hr�8�(�ϲȑ]a��'�QFrמ��|`?b���o���#�ݯ������H�99�0�>��tb�.O@6*�
�B���.(��Z��w�.�m��E�����J�O�����y���������$�ѭF�Ii�@V=�X����sӝ������;�*����/apt�����9t�����0�
E���3{��vS��]���h���f�Q+S-K,�K�I�8�&��&�6�L�6��)�K��Y�b�L[p�^���ݧ�2���%v�G���>�#����'�U�g1��Ġ���'Y���9�˳g(TĻ�p8���w�������Eo�������O�Z���9���w4�D�A����N������Z\^�R�){)�-B���Gٻ�&Μ<KT���g9���ٶ��r�A�h���/�z��G�I,���������Eꕢ.vE',��=��4�JŊ�4��[O�����e'6؇)�n7;wm��}��Ϗ��c���X�y��;O���a�)g���X�T:�����x�x���03�ٓ� |M��5Z�V)���OJ�2_��5`'���
�간������EKKڞ���4*�(��k�L��5�e�{ ���
\�\," q=0:��<�V�.��+����R픍ۊd(o��eE[-���Nj�S;�m��i��0�6'��(#C��܅旋T�6b=}����1k��M�+�f�K$=��0�+k�Q)�k&zb���i���s8�E<�V{]Aa��=��n�믿_@p�}�����_۵0��S��j�t���8��?D�ڥ��2�Z�O?�4s�38=Vz�A�BA�Y���z�����ӛ�E�rk�&�Z�R�J�^$��qV	:��E���	y=4*2 X�����D][�j9Cʪ�5{��w���"ݲ��/��'�Ԁt�Ձ��R���K`7+�����涃�Ь4���J��XO_el|P͔]� ��Ͽ5O>���O�h�h$�E&��f��,]�!v�����tD��<s�]��<a����>>��O*#57}���J뤳8���h	=^-9��eN����S�v��PF!�� �aNݨw���FS�N�q�V�^o�pB������u�T$���
L&ĶŪVC�}�\]Y���նh�de_��It�V#�եH��I)-;]_'���v)�(�o#Ie����ݐ�y(�U���m��;��LDj�#e,!&�m}��Wy�6�6'餔��q��������h�ӰT�	T.)��yu�]M�ץ��M[ٺ}�v4?u����+���iz�c
&��2�ѱd��D��Tf����k+�����e<1�6T�	n�2Lm}��n��@�N����^�N���gd�G��m��),���.kNr�Z�b��;�RN�am�3�r�F݈2����%������S��1Ѯ��窙���}w�t��Tn�Y�$.��/J>���h*y���V�FEc��%�����?�h� �r������s(�Y�R[R.lPm1̖&ɈܣQn�0��K�\5�q��0����or��W�D�Q|n���>�[��Dr�Tv�M[Gi5r�2�v�7����;{���3O�:�8�����8p�mjB���/�O�~�t���t������l.Cu�2g�����<x���l߾K��S'^`u��F�H<�j*�Ȧ[����{LK�tb����x���
d�F�ȧ��q��dT'��(;�Q�HH��2I2�$[vl'><�Z�|6E$짿+D<Ĩ�X�=G�z����n�a��[�*xq�-�f�>e���ա�Zڼש8t ��Ge�D7��G�Ph��xm;�!�Ʈ)���fy�5�൦�0�P*���oo|��K�[�>ZA]���͎�q�UAƋ������D�t<�Q���v�.��9��0���ـ�+J:��\��t"�l���q�"���:��U�&&TGx��e��Zf76W�S�_{o$Yv^�����3k���e�g�,�`b B A��(�bPT��pH��C
ڲ#�vx�a-�B�D��a�����D"@� v�f0���ez���+���V���nU΀���@&9�������|�;��n���0����uܺ7��G(����ζw A�ޚ�cm8���}�ױ9hag��f���8�d
��)l�>�7_����O��f9;
���_x��k�����91n�< ����?�W1I	�x��7��cO�?�i\�~�[8����/|󣷰�:��7p8w�^Y��x���@��wPD*7���b��q�\��ct����$���}hș^ca�%��JgǈʳȢ'��G�
��n�z����q���8:�E#��G&5B-�[�g��O���/�ᦸ��p��&�����-�ֶV1<��J��귏�/����r��3�{�Ү����G.m��p������0X�A�i��bÚ��u�?�����~��o����+-w����{w@��9���7�����h(# �!�9��v�)�F�ȅ�ii1��C�fd���K�tq��i�⹪0���>3S�/C���XQE�f���J�Ms\.�>b(����Q��x������f�K-��:/�^̵)�R���2̨�} ��<��<����!X�l!m|���͆[�օ-����r%;H�=�w�Շ�K    IDAT���zv\ioC��߸���W^�&�����ȅ-�ؚp4NP�:p��u���i��[W������T��u���o��k؈3<{!�ŕ99S��0گ=�<��_~[�|i:���Oa��
"�p�sry)��K�ˤ����,X����bp�9�f�3�||��3�����=O<����w��V���ב�v��s��B�0�ڑ�*�	�uZM���W�%������A_u�Q�';ʰ-����lW:Ўj�$�}A���c8��O�_}��_��W0�{w�_U����4]��{������3x���ɧ?��1���������.�����`�=�������$g[���q��m�#�7s)��]�)XmKS�G�mʳ��11�����?�F+Q[��`~s�g�s��>�%��?�t"��o��m���V����7�O�m�o���T���^z�q�큘�FX��[�R�c�����E������$A��r�0FȖ�&p������ ��A�dx/�՚��@�e51�=��P�˪�x-�Y ��1�D� j-"�[��]�$rS�� �̿X���.������B�Y]��-��T�<��5�k�#m��5J����&������J�N�d�J�D�P�� o�͑Th�v�7�0�60�6q�):�-�?�#A���hx��+��`i�(��x�H0���|�l�I���pxt����[g/"�:�;�O?����<, X�o9
�\��o��9�1�gx�^���_@����������_������/�ԏc��#f�7��_ų�cG;؞�1LX�z^��옾v9��Q�B�0s<���զg4���H�	*ǴUrѐ�.� ��4�E�� ��,�>�S�|��^{�븶}UC9�)E¾�\�}��x���0��:�����(G�+������x嵗��ӏ��(A1��W�����6��y�:gq��ht��g�|WV�������� N��zg����n�xK>�}�9���o`g�>��>��sx��c��L�w0��rLg4`5�#B�3�o�;8��lS�,� �3:�"�#AS�L��
*4#�*�502��l���bI�5S�4ӵ�$��F�+L��BzQEO�D���]�fMa�5�.��y�Ţ��nK�S"CS(k�:�����L�1z+}�w}j��t��� �{�R�/_:�,����;ٿ�l�*j�y$@v<x�J�e�Q���������9d�'#�v'6[��@�%���Q��Ƕ��X��[Le���L���!�R|��ع��x�c-���&ֺS4B󙏽��������tϟ��/����b_�r�������I�^��30�=�6p��1F��:n��U�4J���~��"BOl��`�w�`�7͙lC�z�)͙[o�`H�A�T��L�d+n�9���N�ѳ����)�g���K�l�����dh�'Ù�Y� �t6��QF������îv�v��p�[/k.�J^�8��a�Y�����b��c��34ګp�^y�K�q�sx啯bx0S[��o����d�d���j� ��p}v�9�w�Z�:��s(�s̎5��4�D�b� Š�mD�؏�$}�y\|�H��1��&���Obs�T+9�l�d���~�p��}m�͘��t�q� �nO���ۈZ-�p�d�n�A#�bL�����l�\����ff@$��B1�ژ��aj�.�a�J�XO����T���`�!�'� S�4�6��,ڰ�*�}��\nҶL��u��#'h��W�4������o�:����Eմd��F��BI�#u�|]��<T��q�ְ��;��D�T,83�Uŕ�aM�ټ�:)t�؅�cU"�����!��A����b��%L�6F��ޫ����[�?�Q��}߇�_�qx��/�6v�Z�8���Ξ��h�3׾�[7^�sO?��w����
�|&����x�ѧ��[ ��}������6�x�x(P��/���7��7�]������{�0�x��OH��[�&&�#|�o O�x��#8����\:��}��o!�b81ٱ
���{�y�
�n��G:�g;��zxzuݠ�b�\��l>A�bF�d
s-
;���f�b6��������Kř�D+�U�h�mk��b�yZ����`����b�{�|�7��h�<tD��z�f7�x��Lk���>��>��/��\����Domal�p��-u��ͱ����JO��4rѧ����1�j	|����n�v+Ru�����Vzp��h4[uq#����1�����j��M�g�r����͌�N�4�g�YU�n oF��	9���2U��̙U�������{�;|�/?�k�n�s�&$�T�62�6dC	��i6�P��Qr��%ܼ�wHmDnD����0�CU���u�_����|�� �Gb!]��x�#�}sS`�hǃ���@9[����h_�'�����ΐ�v�l�q<�`k�3��L��}��{�dj��g�Ld�"&�clwƣ)�����K�<�pn���w��sOn rv�'VЉ�+�#r7������+m��{7�~��>�r�����H6,�� ɼ�t4E3l����̾�E!�f��pg�Hլ+����Ϭ���V.b6N�\�Y�Q�T��v�A�!��Q1�3���9��ѝ{�YF�a|�#%��M��6�qVŢ�oY�u�o)ۊ!�t���ʇ�gq8��d/�a4>��,��P��)<۟�(�ސa�CVD��賘%�V���~�S��ҫ�z���^y��4u�}�øw���֦����=�^q��y{U�tr���0��p������akkS��#����I�g���ۀ�/~���y�C�k克yj
)X��^�d`�9��8
�����m5{���'�i|����
�tW��Ϭ=���c����b7=��d4B��^� �W��bL���	��F�&��"�Aę��
������l��y�����Ɔ!�N��s����s�����5�[ ��u�Y�d��Ef�5�l�ʔϘ���;"I�I>� �����k�QL!L��>B� �.�V��!!P�+$0%������8m{J��L�G"#2��b
�;���G�7��[8�8����؏����q���9�7�%��؋�V:^�����0�ǛW^S�q��5$�[8�E������t�>�s/|���/��[��C��/���{哿S���	��`�U��_��Å�/��g1��X���+���}���i��Nw���{��n�c����~��w��=řsV�%�4]<���g�����IBA=���3��\&��G��m`4�a�������M�UŜ�V��]��c��A�f��@���}/�gq���o}M�(���ny�UIϬ5\�����9���<w�4�8�g���a�t��89Y�T����^zY:6�(�H��)YE�o���&#��)䧮��^?>YK�n��G��e��0=��m>ML7�f���4&�6�'��#h��4g��f-�c���S4[�:���q4@�8�1L���1�+mv�I��ja�=VF���c��Yc�� [�/��_��q�Ww�:ݶ
d��T:���읛��'�U���P
;�M���;;��1bEYv(�v(n���&g�*7���}١0�3��`MF�\���4��
�1�h�#��sg���[��+�����2��ۋbO�%���2�F�T.�ȵ�M�c����&C����(��G�[��r��<��.]xR�i��z�n	��6:1���n���b�%�o6��y��Y����A��zp�� ���&�?�f����
>�����4n�c6�IV��v��[��	h�~f�YuVms~�}�-��^
T�J�d��]M~��r���t��Z`7BV�ȝR)̲����\�z~�|��^a�S����k1����� *u��a���u��=b����:6�.��^��h��)q��o~�eܾqk+&�����;�����n$��L�&
n&�)*���H�n�y�vgϞ����'9�V^#B� �G�����d�Ȑ��0S�������&��nl�����D4��ՍUM�X�>���>���^W�7�y2��OP�`^$(
c:M��*���o�R����5pg	u�%z��+��dϩ�=-���N���ݸ����L�b4�� 9����%�*C�q޷0U�K���,-���~��A2��*�]���|�9�_w^�S��f6.�'.Z;T|G@ɽ�p��{LC5o<1��Fj�kkR�&��~�Z��R��<DI��lޒ:�8�cT �v3��"�����Q����g���A��w��	ڃ��@�f���69���}�S�	66�����Ο��+_A�3����CK�H�������?����,G�aG�@�W>���}�w���mƵ�G��~0§>�-\��<.?�D�\����3J�>�s�]2չ���]E��.?�YV�hb������.��R��V����[�K7�d��3kȩ1=$�!��7�Vw%�� ^Q�w��D�s0JSd�&&������^�|���`���xrg.k�<��ߊ�3�㩧.������B�kH#���`p��v��ڽɬ������A���ہ��ё�-r���b^ڠ$S�KL1Lٴ�ɈDR����d�J@n��
[�1��"�M�WԱp��7D�_��c5h� ��vk�%�i�6u2	�c�hl�^A�-)�O�Gc�����O��훶qͶ�M(Dg>��Ĩ��M���ӐQy+���=�H����5�����d,���1y��'�X}΂ ���Q10�=W�^Yw6�x�t�N�R!��OvǠ�2`UgU���G��>�?����H�]�Ȕ'5�dL��g6�p�ԣ�(�2�\D���� �����Ь�m ��z��1;���p��E�����9��Zh�<7ݠ�j���ױ}�k�&W{�Vp<<T�=<��ؖ�TX�F�#G����2��g�0���..^~���H+�z-��_��&��z�g���s��B�5^�A�݃��"�o��'^W2��zs�8��=��]�!׺-�r�j.�P�lk�d���X��zhv���2EOY��"9��x
��E�go����)��w���jsǊ��[�cw���,��R��D���¸�� ��`��-Ǔ4�-�n�&#��#t�!ܿ�GΝ��/
;b���p>�ˎN�=D�J!��h�U���N=F'������TSL�#t�����"���)0+��v��SY9�&��g���`510�t�O�nD��d��cyR�LK���.����Q�!ŷ��񑳣Hm��zd���!5��lf[f
GT�����x.S�,����<�s�#�/6����|:F��})����^�B�����![I#2�,x�*���W���y�!�T#����#������/���J���Yi�`����jꆹVMFc��sO���ڰ�*4Z-�9�.)E�"'l�!Rq8=ƍ{;p�U4{O�`衷z�I.Px��%����w��`�s^���������/�>�~�z������^��}����qsT�I�{�讽�7>���,߷���_��/}�����(v6��
�9��x����x��n������n8�2��
���8�S��j��m�p{�w���j������`��ju��X�^���_�'�KO�w�v0����-	��h=$��(Z&Y�N� S�ʴ@����B�9ܐE*����`�t���l��"�&I�&eh��؛��3�q8q��߾� UsE��Tږ�1ӱ�q����[m �E�b�!�9mF��6�ܸq�t��7��<�;V�8�Ő)R�i�@fk|< d�˴��=�L�_L�Ղ��� �,7.h9B��y2FQ����[Үݺs[ ��p|<�@���8[ԩh%����Vm�\O�� �)�vwU���Đ���p���
�?����<���y����"p���,�FD���ũ�X�	���|���G#�.���rs9�4�3z C���&T!�h�I���K��Vhu�:�������Q{5����766�`�됅 �C%�Dh3��>@��@��*�ZlcUz8�}���pf��{��)ڽ��CU�z!������{\��ޜj�jN�t1X��Ɍ�_	|	�ٳ�Th���<ޤ���B��d�ƒCT��DH J7uv��j��T�����c����Ҥ��.טs�'�J_�\��Е���®�@RDJ���c����{�D��Y29�#l����>8�ֽ=f�6i� ��U�Z�{��Fh5]�y������^��ǞF>�y�#��d|h
�*O��UbZ��У���N���P���A����R����N�3=����`-������nMq�-+#޿�+ͬ�K9��A����w�*q�����ȋ����G�5��U�|��(Z���=] p=J�ם �R��y�<^_Sta����aq_��,.�u"{���[(�&���5u�a�~3r��ԭL�s�G�PƢlq]�\�B�U�t�z����4�d�hMd����%���)LI	�Ě42�cV�@��`71"@t\+����#�\@��Ĝ��Ӥsd�L��& �[�"Z�������:z�A��aZ̰7��`\bu�i�ݝ��	V7�xL?�.~���8.\z��Z�3����V�����8��Ù��{���7���w�"j��}�5<��
��\o��H���0�]�����]��C��/�ѯ|����M��;;K��FO����� ���)�\}��s���XY��p8����jC�T�J�����=�F�p�C��Z"g�Վ���C���D]3f&�u����6~��1^߾����k�6W6�o6���,D��1fqB���L].�ҋ�X�'JÄ���Y��%�+S�셙���#�1�)��]��I�`X�f��׾z�J4�ϣ�\��`h�0��t��vq�j�h��
�1�jA����3m�\����"J-%(�2C#����H��C�m
#��%#hb�Ԕ�,�F�
CBn�6(���*3U��Z�,��;K�h�C<����?�W����?�����Ϫ�ٝ{���5n��P`�eڂXQ�3�;�Ŗx��ߗ��Ƃ�Q�Ň^x?��y7n�P�T2��� Az�&�<V�˯�`�6�5vܠ�t�Y]�H�aoh�~�.�q(=��ޣ�c�;�#S�|�H2�jg�����='E�
nB���@�+�	 �㑩��Z��uc��n1G�ȴn�v+
.�%��dS
D~����*S�3� ���_��g6|��kOI�v�L������(���1�aG��,����R7k飜E�
/E��*�.+�ٟ�]!x�{ ������JQ*���@`	7#{DqFҒ����TIY̔����D��C�t���Tih�ژ�]��}�hG}M���khv|d��0�N��D]NȠ��u/$Y�3[�`{g��_�"��̆8�����}��\׎ � +h�0gQ�E�Y���38�v��ҫ�{x�����#U)�?�G��"�Z�*��m�'x!����&�)mV\�d�1B�M|��70�"����d6�x�=�(fC�n��=�1r��|p�F���]�������
�{4���͍n��>�f���0]j�KE��D
�\��0)F�k�*���y��7�����>�s�l���>���.����FR��=���Z��Щ���0��C$Y�1���@a�������$y������,F���6��I��~�4Q��x��7���/������ �=�&� 1[���M�;��\J��T�Z+5�����`<½�!:+�Pz}ܼ=D���(� /]������&:�˘���"��əu��}K���������m�n��w���c��#��Gb	��YP����Ͻ�ѥ��]����7?(������n|�7|��lU�zu�N��鴱��'�u�H��q�(�c��y\�rM�@o�VTٍ}w�S�6�ٗ�    IDATO1h�*�44��C��ag�V������,qc�^{�����i���2�=3���f����%�h7{Tr)w�K��C��ϦF4��/�H��hw���,i.J��Zș�LP�:1/1OC���m�qm�����&�d&m����|J�5��R���(�gO\c��Va��~a;9.8�rS4.�,^1�0���~���U�S��L�Ux��)�.Ԗ���*����'�p���LS(��t:����.��;8������ƥ�^���K����F{��:����\�}-���+����-�F��z?jb4���*u{\�^~e���U����������k��o�����><2V�ɃL�i�E��x<F�nu��z�1mƔ5�J��a4eʾ���U�bc31��X�Gv4K��~��jH2�>-q�G�}`ٗ��!Y�&���4Ip�����J����o�=�X$Pe�5}xE��]t.z��N�"�cu�A��K�����^����"ü��dC�ޒ�8�&�ŹM��7$ìJϜ:2c��7[��s����Z��+b�D���J�q�&/�T���:�@)b���r�9ϔ����L_-&�l֮�l����8��A��c��7��a���@��[:���IQ`������D�&s�y�N���g�Ïy9�����;{�jm� �6[x���u����pv�^{�%����=l���;)��n�m��ҏ��[��_�0�F��G�Fs�ߛ��{�4��=l�u��E������64'0�i
��ja��l�P��lz�fo_�ra{�_|�~�88z/|�	�ľ#�SQ�1��yU�j�L(�G\�X,��Hr;�	vFZ�~��E[��F@�����
�?.B�A�\s�؄�%FZ��/���=�o��M�a�>��b�xٜ��^]Y�f�'���Ą��ua���ۻ���?�|^�Ν�i�T��	DX  ���,k8?iUU���
�8�׿�*��>.\���"��z�	x��Lh�ĵ�7`��IZ�X��5�3k��D
��nql+JRX����>8��h���9��:�lq��S*�|���66�#�P+T�Q�r��|�~O?y	��p�������!��i����E��+/��|����q\�<�w1
���_����O����m��-/LG� ���Nw���1ಧl�7��`2	pv��m!ƭ햇n\"φ@��ۧ(?C�L�,� �ճ������֭֘���^�\�*�~GS�)�M34����%����&�86=r�Y�d^
%#�fTM��0%� L!W34��R\1ө�3��w�
�t>+�-CvdpZ�W�㗯�(6ά��{b�����.��Nc�(b��D����5b2�F[�bi�M*��i�ރ��Z���J)����X8:��\m�}̦S�0��qb@S+��Y:{���8n"lrOƐ�y2R���Z�^O��	 �q��M���F��[����*��.\j\Ly>��=�L�j7@Q�g��/�� �<A�'����#�{]�~kWm����)٬��l�*�)�y�R�Xg�#k@��"� ���-<��1K�dŀV��㬠�Ӣd����<���M����h��2��pj�?���~�����:�qVX[oc�ґ7�ʠ��EQN��4�6� Z���������c���F+^>���.:�>�*@1+�UL�2�Ů
�$U@]5x��.�U��yE�p�����*#�&�H^�s�^��Z���Mg�'7q�D#ħ��t�8�k���H�K�M�IJ�(ZM�}2�'�g��J6�����L��j�%Ci��d�wzJ�H�:K����dʤB�_��l�$d]��z�5P�)�h�ȝ{�#4{�� �0�Ј��N��tq�(�Q$�	ШG�xh7��@��c�[�62i�2�A.�t}L�%��e�/�Ё�a�EF��:�F���.�xI�;�!���+�*6)l�q���"�7o+X���h��g�XclT���3�1�(X��4�1&��i�b.cfW�`안�����䌱L���eg2d)q�����Q�o��&��X]�!�l��"p�)Ƥqe�R�R`@��0�R�w0@�Y%�p�xl��#�k+Ҝ?,�"(�uk�V�upc-edg� �qpD	
[�N&���,{�o���
|�TH�Lu���4r�9�4R��)u�dU>����A��!��<����!�.����x�y�|�?�k7�˚�!���m�~����,�Go�	v�i\Mh�=�!P�|�o|����RS�.@���[
~�3��[7?�뾿�ƴH���196=n'���p��Sx�k8>`C�0X�c�՘�=�������9|U��`��p���'�@�_�ʹ������4b������5�h�[��cT4��&p�x�h1F���P��S�,�D_�l�K�6{��h��QL�2E@��=(}K=�V9J�0��������8g�G�O(���{4���lj*b3QZ4�.��a*Zm��"�t�8���i6�~��4S��$�#2����a���0��S横��@S�&�-�+Y���,R0�����5F��K��
��x�k45U���<�d,� �F���h��"�(:WQ�9S�8mE��*����dz�v�6	\V��}�6n��~�6(mi i_3:b�_�vks�Rt.EQ�;�(7ۆ��&��VHs2�9��1�s,�fӑ�.
C��4�&�(�`q3��Ȅ��M7е%0��`���i�Y8Y�7���l�/�d��sz��&�*C;r�Ҏq�L�K�
�Z1B�C��7��!��=@�d�'���]QQC��CS��$�u�����b�!�=�ې-��7p�n�9%����P�SsS21~e�1!0V{3���L_c��]Nu��4�dk�b+�h��OPy���Z���dh��,�����L�g%�C$�	���������S�9K�Q�ud�JoE)JVg{d]w �Ȁ�Fp����ך�Okp��}L�R���Ӽ���|t�*����5fdЀ���|�A�����,�#��������v�c�?=���1f�8�q�͊m��ҹ�Ȇ��o��tUe���pp4�����ҹ3�V�S�A�+�Й����ӝ�*�K��#��a\8aQ�#K�Y2�Sd',&�֦ٶ�3f���b:]Ef]1.\~W���������@�b>��zg
�M!��W��a���#ӭ�~���KFHf�ٓ0�ѻV%0��5t5,��2id�Yɞ���j�/i�s��ڔS$�Q��$��dI�m>ݸ�������Q�
��	����S;��dU��k�����m<�)q�̓���5a�����;���A�Np��x�����?�"��z��2<@��ೝ� �Ȥ�E{����������?�<(�����߾���p�����c8e��l*�ި{;����t��c��HB}V���5QO�, !h��&If�qS���Z��e2@��p#�X���񢍂K:��a��c)P,0�4�?�������ٰ\A�)B�_��r�g3tY��J�F6���(B�:jPh����[��'d�2��X��
8�3��2��a�d�IO-y��ki�J�Z�̴�x8�L���bcc��:23ճ`&1:E�#�95����t
L �*�g�Iy�4�f�Jv�l[K��&X�G`e4�|����\$�ip��{�Ԡ:��`�Ѷ��у�@�c��ۘ�ڤz,�A	ܥ�$�D:Ќ#�M�d�ئKV4��f�se��Iѳ���!�@�R,�j[O��$p��- -Y98|Y���D�y�9v�@hF������i��`��+�n)��`�˔P�Ȃ2� �ҩϬ˱���\�@��;2y��|T�6�@��IƜ��J�˱�ZE�g�96�oێٿi^���i������o!����9-Ω���bljo9��2�Ӈ�2Ӣ�hQ?%�X�W��5����'1��S+�Zq>F�H�|z�1�o�N�-��Z�U�����ԛ���)��vo���j��h"[l�����O͎e�,�#�G��0��fH���9�>�@�ds�6�	�Pf�s����Vq�0���<���Ɨ�F�����qPkJI	ǘ���\�����2�A�̭��\;��yb�<yӳ@��{�F�z �2���KZ鹺��ǃ�w�N뚷u@6�4'�����:Qw%��r���z�u$;m�'&�n�i�i��l�Im-�yv2����}L0C����m����]���y׽��;�����z���cA����������p��X�D�b�nKa�����}k�JNf贺�9c恵�gx��h5=�߾���}�l�a>c�L^�ͷ�5���������C��;��G�@�׿������~�u�>�ٓ2gk4ڶ�_�+�������Y��&m3MvV�
CWv\�bF�ә�a?>� �S�~ˋ����Q~Y�Z|c�3U�Q���/�KKmM	�f�S�%mB�,�;q�H�������I�MW�%˄d2CJf,�֌���&Si�j�dBM7CI����a�LYV�l*���B	d�������&ө��ix^����V4i�v�&f�����5��N(uTm6���j �&�w��4�㿹���~Np�zz��͢��&�h6d�8��`�6�n	���~ou&�"���O֔@Il!;;�c77�L˴ �jF�	���(���U�xs`�|I`�9DƨІk� ��I{(0i��>�f�\R�I�Am�B�ܳ�]��9���:8C�԰�d{fb	�8��G��C����n5�F.3rFH(���o:p0ZR������=3��9|z���Q�B4R_�?iQ�G����S� ��0mz��y��Y�O�d��^3c�4� �mkf4�F�`@�}�T��)�������c=�;m
��Î�iG�(].�-�A� T�:�0(c�����2��dz	>x}2���F�0҄��d�\������u���C��S�z�jy���.+�Kk�٥-��f(���9a5�R�������G�q�>����
�B�9����S5w���L (�k��,�0A���R'�U�;2����xR"T�Z���<U���	�޾��´����yc�F3���=���H]x�	ۂ2]+����vg����TxH=<ǟkK�ili�욵B�ǡ&tlu��6�d����Wr��!�'#�ҩ
�$�(� Mk-��*n\��8lI�þ����^�6��0f1��c��R�*�i{�k���s��.ͫ�בݻ8���_��/�������A�SQΥ���*�7W]��Γ�*1iػ�[�
�`����\t��#������b-���aIm������̅=�@&I�-�X���$`:������=?[i	.(\pX%H����;7���Ȧ%U���E��"�l�:� P�qA��Ң�lR��A,��|¢�b��Kf�V�ʈ�58�}C녗�B��,+<i��BF�jq���CqL�1�;��+f+��ip��f���Y����u;)�0���SZ\��'��XȔ��bO�F��ݨm��Kj�mU��;y��o�.�f��~s�3�x����
�ӡ� ��C�K�%_�S�M�n@,� �D��)N�ϢF�@�>f��R�2�����Y�L?Y���f�ͣq��CQW�y�b�i�2�u�~�6�s��*q��f��k4h�A����&�hnW�)�4"��L����y�ۀ�E��;W
^3~��>v3^�d�5�\ۖ�׉�S/���i���͞zBJ�O�
yM���:ʘR����&h3�an	D���5F��E7ƾɎ��O���3:R�����l'd��ap�v�U�:��T���� ���)����"�%($@9���,���q+����s`�W3aZ,���Q�����|����F��3�/6��R5��U=��f^3�A�.͆�e��.���d�9^�N$	����j����35���bP�5��3�Q��wC;m�c�@�m'i[�����R<NM��]Om`*+���VA���gh5LF����^2�5{�`����P,dLɑ��C�Mk0��,4cTF8w'q*�"AAK(�7��߬��1���!-Te��dCC�8ґ�����n:NА�5d� A��ŋ���.0����#�P��_��x��g�ϸ1�OP�4NE7�<�|>0��7� P�b�svu!Ӈ��0��i�J���cd6K�d�#�7rÀ(�bP�W!��q�+��)nPQ����icX��QV�%�ѸݴN�x�E�n|�93	�-3�M�7SHB�j���GSg���0�6�����FŶO�]��F��Qb攪0���-kX����|��*�e�Z���zA�yJ�Znu�P1,�l$�sL�#GN�,�`%��
��c�_�̳qc2e���_L��,s�F<'�:�S�D�R�\`��D�����i�Ǎ�fp��Ym{S��HU3c�O�Y=�-��Ӭ}�TlC0r�3��L'2�+fh����54E�Ɯox<;>�
G�g榙�Ɨ��6r��6���u6�� ��O<I_�{�'&�2C&�#��l����P��Rm�,�7e_Q�XϨ�`�l��^�Ŕ�⚨���H]�i�v��Y6�)�xD�10ޗ�{N�=uq�`�߃�6s�a}Mg<������o1,�O`X��J�s�İ�E�`�N�r^��`X]n3G�b�C��Z�k��/ٰȩ�ʰG$Y�ւ��-S��k�cH+Xs*M�d��]���Y�\;�p�-�c����SOຣ����=|���V�A򆪵������U���R�Z/صĀ-�7���@]����`�3�}��f�,��f����m6휳k��v��5ð����75�T�AV^l�h^��f�o|ތ����Z�f͡��/c�����Q��"��H~����(��b
u���{%�\��#S��u:U�hf1̸U>�y1����&(d���0/���;����K�a�C/�#��޴#���	��o?���;Q�������#�P��k_�g��۟�_[͹�I�G{
�e���	��H�mDs��$(aOv�7�2MF��hX�X�T,m"\8E��$��&gj�Di��M'F�2U���vv�5��ܸv4��W�K�)���E���6�zC��H�*��FO���G�Iw����dL5�IC���\V�Յ��u��X�F����1��c��^���,�i�ײ����L�5&��p��ZG��l�^,.�'��6I;�v��1F�P:�:����4A�L��Y�L��ȱ�b [SYivh�R/�/��cÖw�z�:;�G ����T�`�\��ޖ_�UL,x�8r<�&4)'V��R&8b^���P���$�����b��86-	�j)����S/t1'[B�8����y�(��x�X'�$cy�ւ�L��6>�2φ���BPh�c�ӯV3h�� �`7m���ȿ/26�4��3i�S"���b�kl{����~���Ђ?��	O@�C�Ƕyd{�.n<G��9�j���M�`\�8�:Ǧ-�h��X ۿ��4:�A����v��\^dL-x:a�X��Sz�>?����F��ڵ�+��ƺ���{�t$:�;�9g�Q�C�~����H�h���!�n�)����x��#(d�c�h�����n��~� �?y�����������\�߹6�8,�K2;��Wd���z���oE�I���^��`�VE���f\�N
{]8�W�jJ�d	zbJ�Nm2ׄZ���1�)��4ǸL$�����o<7�3�o�d@'��5���=�A�x�����m�����B���`����x(P���������~���I��d��We� ˧�=���dZ�D�v��)fﴑpq�~��*��B�!+�V����Y
��o�.�1���	z��p�_�1hV3*T'��j�����Tk�qqA�`Ħ��a�J�������̱��g��� 3����^����	��sJ�2��>E�5�MB�]�N���� A�+�âO��  �IDAT.j�c$O-c�ɘs2)�����{�v�\�T��9����-i+��"�T�#� ;ضt�/�,שIvy�d(2L�:���I���!��@�_���C4���Dыj�������nY�E��j�[l6/�_�����ֆ�����Sm<�,�%ȴY�#��j��
�����w�s
M�kM���*R��.�w�ˬ�����Pn���TQ�:�����*�i���,��ϓ�W�G�%���n�g���S@��ǵ�)[ �0��<�~�>��a�S�+�I/j{m:�)x++!��)T`�4�!M�Fтc�S^�Լ��҈��cXl�U�O'�|�	���.����Xh�ۂi�X.Sk�I���[f5�j6�p�6p�p0�7��+���i�f�)Ku�`
��Z2�%8d��I#�Ըި�_����O�~�#i��>g nd���DEn�
Rk-�)P���A��Ź���8X���\׾f�t���7�&׌�`�������)Qc�����w�����={-,@�.��6�(%L1Y�X�f/�3�]-��^a�1-e���<ǔVX�#�%<��ǌ�����͏�W���������i��{�,O��F�@�������7~�ݘE���r2KiE3E���V"�MO���S�}�T `t6��MJ�mF�j_L	����2�]�Y1Q�*5}l�N0Hވ���djOf̛i\L�`75�[�����-;`��ԝ���pq��)�H�I�cV�Yܡ4��ޠ���v$�B�ة��,��?�)���16iV��zIY��o6"k�W���bA�m�ٞ�='�ؚ�ͤ��w��_�^'��V4�ty�60�d�� S�p&Ǥ���1�`�0�`��|?S�\�����O�t�l�� L:�Bx~���0Z��3d�ޭә$0�O�d
F,�y�������0�6 �R�иupR�r��Ƈ}t-cwzFDP��l�FE���,pX3��a[0��0%�q�l�*fS�$�a�yk�m��&�kkeqN�O�
��V�y�"(���<(ٚ����攭9��?ݐO@��A�)�XL7����,����T��uJ��ީ=1-�R���#�m��n�U���{�W�A%¥UE0��>���w��v�5�TmZ�`�bx�L��9����;Y0�G�9'� CO���Q�a����4�s�g��H�<���KV�x�����Sp'�N�v�fjpl�L��\7u�mx\?�`v�l�{/�y��~�X-5���ׅ;6�b|x�`�q����7�U��|o�O���6��m�!��-0����^SY�dF�@�{Г1�����2G�30��^�h��y��WʫU Rn
$0�ZIK)��]_�$���?��n���'�m�1��r��#�P��3���?���ʯ��dӭ��cIV#����uSu8�j��暊��v�75���ѕ��<���I���!�c-@�� P�ݏ�bd��9Fo"sVm��6����3�#�$H�BJ6B��I���� gaI����uz���MC�de�y�	2�O۹��NOфtF;��Y��㵬��-�i�g7���A�!�l�uTq������0 ~�~���luqҨ�
{��&B���6Ҳ���D�Z��C�� �F�[k�����96[+֑f�v�D�㺪�ce���1sH ��Zi�S����,��]a_g����H��1L�I��m�����\��Y�`#��N74�m }�����`L;��y~R�C��r�.0T�	/j�ئ��f�~5(���f������������]eu�w�^d������L퇧�Z�1�y����cY5���X��w�E����Ӡ�0�6p���f�S��`�4{�8�-�h����G�jnzu/��Z�kd�n��NPk������.�-6zJ[c���k�RQ�X;��ޡ����0S���t�0�7j��p�L5{2�d�jfͮ�բ���5�g���q���0��2�����]���#S`#�Tzk���4/-vנw�j�s��e[�}A�
f�]Ԉ/�*��N��Vx���B>l
>S�W�6�+�Y3-ȷl8�A2������:5�T�e�e��p��D<>�i��&����C9��`�zh��9�JO�����I
����c���_����?��Ϙ*��c9�x(P������|���c;��Ydî��b5�����q��u\%��:NU�6�Y����fVU���8\_���D��\�)X�%	���R䍪���Q��*i�U��-ۊH^��|]�a�{�SjE�I�N���H�;�W�P*����%��\O� r��)���'![V�NV�.;mQDY*}�gy��S�P9['8�Cf�ǜ~��-\�-9DEQxEQ8��;dѸ ��,c�yn�y~唬9��3K�t�.HCX��λ,u:��x��	�����]��H�m<ʢt�ԩ��kXY�n�hWEQ���U�c����s���Z�J���R}7*�N���F���7Ͳ,�$I\�0��s�0 ���pX�ᗥ�j��eִ�Iݑ}ʩ�G��s|X�NX������Vu���[M������Qƴ2u��5`R9O�� �S��9�����w̘�߈*6`�2��,f�7x��X�#����{O��E{�l'S'��޵u7��}�0ԧ63�~�FTJ�T�0���MV���Z����\/�"i肋��"�
z3�-h����@��>�-���m�j�-{tyj��"���q谍f�?M��Xhc�E���T�yH��-�a|��w��Y�a��	(�A����fQ��:��{O�j�I�/��ebi4�*�XxCi늠���M��S��e��~�"ش�WkaC?�E6Ў�a?M0���"h��Ԛ����A�kg�(X��#���(=.�^�s��u�F�I�۹o��k��<?���X`o��
���BA?�ej�G���P�%k0����Xw ��	^kͮ��5i�zU�<���>��>�}O��2}��DB˗���C�B��7����￧z-��#��c�t%NUH�a�<M�W����B�vU�,]�rK7�f��W3ߋRǩ�ҭ��tܲd���7P�|��
��GH�q�9-���x����N���s�d�X�)��g0�9G��NU�l��"�Y\�:A����<�*�*'F-\����0�m�<�/����ʯ�jV����%�ps�ȝ�^_Un{n�zEE?ל�ܛ睠U�s<��(湛�3��|c�4͙�+�fX���y�8n�dy�UeY9�9F��l�*t�|V�e��.iA=��|[幮�W^Y�L8«�p+�f��������4;l	��T�	N�N�:�!!�W�e@`�W��9�O0��(K/��FQ�nE#G��dQ��k�:e�y����e�g�+�T�eQ�5x%鐗���K�XP4£V=��L���B��{����́�������V�hF��(YRpzI��a�
��r���]λ�ϗD�e����v#��iS���q\�����}
���W�E��
iT��@��*����æ����y`�I�����]VF�n5������2dT�M��y���X�%wY�?}e �����Mt0:
�,ʸ*ʰ�*����*'/����2�=�QU�EjH��[|��rY���][*�L�Xe�7�f�_��MNL���gI򍤋�#�E�RF��.e�zn�:l�bⰲ(8+N%��ȭ��I;*��'�]�v.<iK���#[syp1�*2�I�/^(��^n��̓����??]�Q�3OfF|l@1�R�#a��fݎH�:=E�|�$��(�Ǎ����B��TU�Βĥ4�s|�t�$���V����~H��׫6ou~??;�R��~�"e~t�p��@��J��+b(���êo�-y�y�ȌU���K������i�S� ���<��W��t��|��ݰ�:�r4��|��3��1TSV�P,lDD��ײ�`�nU��?�(KW+P��¹V1��#,��W���j$"�'v��e�����Ne��
�����sq�@inx>�_�"�f#�s:)��Y�)�Х(�</�"�4^^�Ճ�R>���gLt�z�Vi�������ZPNgL����ow�����O��g9;
���[��r�s�I�����o�㿟q��>�kv���V���;��u��\w}W�������5��>ww����*�����e���g \�N���������j�*˴rwY
����y��������{��^e����,ϋ+���R�㎝�l�䎝Å!��,��Za�j ���3�;�8e�U�˴:��㺡�����*�{���w��gU�>йs|vw�(��y��A��9N<=ߏ�ĵ��F:'~�ƦL�k��k\��Q�*�gz��(�\����s��9�p=����`��4ϛ�Л8����p��ߧ1N�$)�v�1��ơß|mQ4���~�Y����������7s�<���xE�Qyc{|���ׯ�PϏ�>_k�k�=c��|�! ~����9���%כ;�8^b�r=L���=�$p8�\/p�Ɍ���Q�@�������S��A�ƄUY�Uш*��h5#q�z3�ug�� ��g�>��^ߎ�v�VeѨF^�t��A�kU���â�UyީVV�2�'�[o]��~�ї����X��w1x˷.G`9�X��r�#���X���+�<��,G`9�X��r�#�.F`	
���-ߺ��,G`9�X��r�[F`	
�[���<�#���,G`9�X����%(|��|�r�#���,G`9��n�%(�n����X��r�#���,G`9�b���]���X��r�#���,G�e����J.�c9�X��r�#�����X��w1x˷.G`9�X��r�#���X���+�<��,G`9�X��r�#�.F`	
���-ߺ��,G`9�X��r�[F��c��(^KV    IEND�B`�PK
     ��/Z��5�) ) /   images/fbc1041b-f35a-4c82-8c92-5608856c8a22.png�PNG

   IHDR  �     ��?   	pHYs  �  ��+  ��IDATx��Y�fi����ߗ�##r�ʪ�Z���g�3=x��!\�� �����Ȁ��H !.,@�XF�a���i��{m]��UY�V����������#s�c	�}���PDF����|߻<��������������c
Wc5Vc5Vc5Vc5Vc
Wc5Vc5Vc5Vc5Vc
Wc5Vc5Vc5Vc5VCV�p5Vc5Vc5Vc5Vc5d
Wc5Vc5Vc5Vc5VCV�p5Vc5Vc5Vc5Vc5d
Wc5Vc5Vc5Vc5VCV�p5Vc5Vc5Vc5Vc5d
Wc5Vc5Vc5Vc5VCV�p5Vc5Vc5Vc5Vc5�_(,��y苌����5~׷E������g~��r��o�R|��?���]|�/��|�3�ӷ^�2~�����2s��xq�+~>��Zn~���.r�����g��#������#~�˅���ef^�����/߫���c|o⫊�������y^X�_��Y��g�����y���6�w^~a�o����c�64�����y�r�HG������_�AI���h���=H����g��jI����~��_�yIϖ�-��Ϻ����|��\�}矞�[/փ�[��߿��4���e-�|��_��e/�P��WC���/d�;/d�R/e0�
4��̖[����+�@b>�zr�gj۶o��~:�nQdE��_\<v6�J&��Y�s�0��"uꍆ,��3���従U7˫��Skf[b9��m��ȩI���Bka9I�FqjGvb5�-�%ka�/�U-�'�ٲ"+Ic/��/�"�ݜ�/�z
W.$I�-���
�xx��ev��4���d�X�׮�����ƿ��/
=��_��}������kg���D�f}fY�7�ϛ�� Zǲ�\�GQd���
�>w��^>�k.���T+�i�R�tŋ�l:�ǝf�cU��7M* |kkk'�m��}�r�Y�&�}V��^����ĳm/�<+�1۱��l�%���[��!�eR�����Į�F`�<K�,MSY$��1�����q�aJ	��ˏ���R���N���j ��v��OjA���E{#��8���UX��y6'`a�E�ۂ�9?�������0�;~��G�����)���O�k/��J�dA�gV��Hib͆��x>��j�q{}c�XE���3�<O���~�����kX������f���~�9�En�Y�|�ӿ�ʙR��3���|>��_�p^�[X��*���iIͯ�O?�ݘ���؉3�w�d�k%zYƙcb���d���x{� ����:�w|.�/�u��xbb�q���x��d�����' ���ųp��«�m����WH������b�k�ܙGa5�� *9^��i�s �Y�tceI�Eq����v02�sI>.֢�@�aw�R���������"�+��7�z�X���Q-M��� ����slr�?2�H��r9?�W;==���t��c�񰾾�v����E���>�F�����r E�8Wt>X<��7����E�Q�1C���xN[��f�����a9���[�J	DNu��������ϙ����<�,���7��k�J��������|:md\[�<7���I��ꑞ@3��$agy�z�hQŒ��-0!|�?�o�=ߧ���N�$n�f`U��ւy�����0�q@�n-|e�<�䜟�*9���Ե�k��d*I��9�@7⺐!.HtF����~լ�e�+mP���T �%��I�fY b���^
��Xk@ݜ�
�3�T�b2��i�ؐ	q%�sN�BH���{K��TV�BP$�3��ż�V���	L_���Nb����jB@������y�=�;���Z9���i���������'�MFPT
༔��Y�w�"dn�E��?`]�m��}mn�����$N*�u>���b�,�����~��������b���o������Ł�)�@������l���>/l�n?_��5,�;	{q�Ԯ]�~tvv��_	��y�|ؼq�ֳǟ]4IǶ�ީ;����s��,㺋0����h)^Ҕ��ڤ]hK�%�u�@ĩI��]|b ��12E �#ʫ6d��߀@��E��{��l�C�C\�h�%K��ET��<Ļ���"ZȬ��;��?x�����x?y뭿2��X�W�
?�࿽���O�fŝ�k���S%��BIcG�N���'	9�V�)�V@0�4�d6�b���w]�$�0��d�xҗz�*Xk�@������ٗF����g�>�pK��|*��lI�OUE C������߫`����`X}�8!��X�!j埓$�9�8�-��RB�&J���"x�P�}i��Y9�01Ap���s����@�X"Mc�	
��B�Wp��P���y������`,�VC*��ηw��<.�=�,)ߍ��+��x<�<�63�1N��bQ���-���ҁ��ޚ���Z���$�}�2�$B0����I�0�mc�C�
� �yj�|m��ˣĢ�#cօs#dɩ�t�9?@�(8��`4S���N����:Y���ӦF��\��,��o�k5�8^e�kϵ�w��kC����~��C(P�����b���-��πI��<���t]G���q�@���*N��G�(�p����#�A�M���]��,,��g���>���{/��S�"��h��{�{� ���s�9�%���X���N���������~||��,�V�Z+ �0'>�	#��P���uyy��M���#�>�`� ��źX���Q�.�V�9���s%�p����
�j@@%B6YD>�4�>$��B�z��^+ȱ�|[>�I�T����U}^B�V~R��Jz ��sj_�g���� mE����Ʃ����!_<��㞀_ ΄�V������M�Y��X��<����2^���<��x�=��A�ϣpn�������cd�C�p���ˍG4/�-T~�{�����si0+�����9�IC�fS�r���򽮿#�D���.崔2|)����J�ˆW0`)���~�����j�*������Ǻ6��@�4���Mi�+�s�m(W�\� ks|�TiH��PZ�s۸����щMs31�x٭m�_zM��:�T�q޼W�� 0�y��\�E"n�
}�O$꫹�T�,�.DnL~��є�F[�?}�+����p���|-����?Psv5V��+��(:�����v;��'�JWZ5|&���h���ݚ�¹����d<J���Ϗ�p�<�J��U Čd
�i7�  �-"iշ��7ޒ(���lr �(���J���f�0F��fr�#�t�T
e[(�N`��9 ��"+ <=2�R0��9U0�eA)8�.��|��C�N���Ršߛ�L&*�����]@����,��A��U&(�R潨��[����L=X c(�*�T%��78xO�l�
������ߡ�-_M�$���6`��'*h.+��R0V(��u���VG��Βԅ� p��nL��(��(8t��(�T��ؙ+K��Q���/�e	P�AF�)l�N����a��`ͳ��/8�Z#��F�}�3s]c+S�>�{���R	)���,�\ݒ��P�Rz}f��Tl�Z��%I�e#^�R��=�2SZ�^�ɯk�{��뽶��R*H*y	����Pú�P,@Ζ���4l�!(�V���M�]!����X��J�-�,!ȴ/�Hj��<����I�Y�(d
y  T�-���[T%���K�֔�td֤���/���q$ ��e8
2�̱�u�'�� �H��wl����
2�  ­�����N���+��!�kSC��� ;��B�/�K �.tY��AY����z��t��)�s� 2����$Q��|]��Q��.����p��d�02*ɕ�-��o:C�G�Հ%��`��׵�� �l�����8�5�
�����)���3�oj��l")�4 ��#���i�u N�� ��"�󰆠��`,^����U(أ�,��a2c|p?�O���f�r}1W�V0A�= ����	b9ϐ:
k��&�$x�f�!�ۻ2O)=��詜�ci7+����>�����CWŠ�J)��r�T�\�A�t6��aY/����1�uO-W� ���Aq�HLP������-��j�x��4\���|�����@�U�At�?��Qm�6� �8��X�W�
7ۨxV+�5�٩"��p�J�Of�����US��r#�Vu)]\\�ث�_�����q�֣��PR.�-s2`�5�m����>>ȝi[f�&��@��/�	�B6��~G��5�s&�V�M��Y��N��9�	�h�yP� ��G� �ʉ���j�'FU��
�JP��ʄ«UTp�l���/�/�Uf�,H���#,�k�1 ��n�x4��xȿ��^��0Q��Ux���F^�xRL�v_^(�4�p�B����+A2�a�%ƚ'=aܬ�V�^zzx�f����K��/��R�ӻT H-���S�@�b��~iMD-x(ǀ���T=���!e:�j�C���	q@{�W�ҭ���� ��$S���� {SҴQ���� y�9�#��n��'/�}�P-�$�+W���lЍ$�ͥz�	ְζ�25l���GS1���_ߗ������]y��Y__�w�Mf"��k�g��z	j�$-���z[y�t<�M%������k�%���B�}y�3Ҧ�5�����QB��F�t�Q�نn�ңEPz �� �C��x:��:1�׆�����v�ٟ�����SU�|����Z|_�=R����.��� y	"�.=T
0i<�yΟ�����ť�d<�/��@~�����G�~$�+ޏ� ߕ��@��ihɗ��咦�W��ϧ�wUl�s^��\�+��z�5p�=��VEH�r=����\Zz�U(��7F��>k� }�z���n��ktv�Ht7��/���ԕ��dv��U����/�i�ya�X�m��K�B>w�f^�/�t����#��/z���#7��!�'}��}�M � 4�ej<���%廛�����K��Kr�Ŝ^����ҋ���|_F(�S׬g@:��/|�f_�ʮ��X#��_���F&���2>;���6x;���̝-�w7��\�(\�W�
�Ԯg�ȳ[Y��-i�6e�*���|�p��r� d-yt�H�oޒZА$3%MiTץѓ���;�e�CYN2��Sۖ�,��{����,BX��|�l���	O�22�Ǭ##�,ep�zs���O#���0���g�؋fz-[��1�[�K P0�,RO�f�QH�x~�Тm�POM 0�<%�W��b��SWA�o��(@6 �!Oꐄ���Ԛ�kU����s �f�"�F� z�J�HO���P�`�QJa:Q�ݯ��ԗ)�����𞫾&���D9����GeP���2�[U���|���I`a6'#���:e�B!��t��>	="t�f�T�R��
�ԃД1��*=�Q��~MAh-�.I��Sk��F0
4|���u�Kţ
k�����hQz�l�"U��w!h�S�R($�q�E��
L�T���I(7v�JÁ�A�����vϰ�㹾/3�< �8��w���;(�aN��+s"�6���H�k3G_�Y[�rnB�^�sSC����/cxq�k�-&�I����<|VCT���T^�'�?Ґ�eN��ʥ�K�/He:�k�#�w���Mf㑃R�q���\�ih��
�I?���Oa��P�$��d%O�(��-5�OS�Fciz������i�p$o������-�mF���w(\Җ�`TA�*u#����~tO魧��"H`�[ԛE��i%j�� �z��w�� ��
���(V �C~XP�I�#���e�I��K����Xee���$��
c��G���_�s��` -��o���tV������YL�P�!/�& ��4���ꪬ[��X�u����	�\�l�� }�?�ノ��o����6��k�`��Kܓi�d�{$��,|n�Ɲ��%׀���4�Ť`m3[=�v��G�����d��辳sCl��<�|*���2�cy�krs�"�uȱ��ЕF����;eS7
7H�4:�'�p����j]�8Qc�,�f-��-$q}����-4��ȵt�d>Q٥��ܔN���9��dd<����k����H��?��n\plKo:��Ɂ�oMR��5�\��)�DVc5^a�2(�����j�'��\��
� ����-�+M9x~l,'0��{M�|t!���ʍ�+��\�;wߒ'G������{&k��lt��Fy����	+�����D=8��>�����2��lkޔG�"Sn��\\m0QX��l#�*]�w�v��)AK��$a�-T��������w1YH�6^
(좪�CA)$׈R=UK҃B�͍��p�Iv�J#UVih�0x3�g�	֯	�1c�`���aO@+n��C�GP�#�4l�!J`���'��u��6O�9��%�Z��V�����,�4�T d�S
�`� t:�+�����榥 ^��p0WM-g[C8�+(^��l�YW����	s����E��H�f�=NAW�[Zkt���x��h��V=_ n�^X�4O˰����8����V��0�_0\��h��PQ���[z��t�c�{hXH=�����b�����B�0�:�z
�X+	`�gQ��K/�����	�=�����2.�_c��G	���0-!�"ϱ�~���w���-/  ���Y@�1�k��\�|7��2Ae�`U�����Y�^!�뤯�0�쥧��U
E�gS��k
�
 �*��&�)���6�-� `Ӝc���J�Cp�4�6��b��g3]�aS��&X�����A�зO��#��¹��x�YK�$�^�����һ��wۼ#Y���LZ�)2���˥7�R�&"&9�� ��S;`,����<q�$h�D3�uQ*��9p�����^��s͗� �-+f"@U|O�� ��>���e�����yf�蹆�-Me��R����B=��a��Ilr�	��[�bCe��L���$�XsRz�Vjd�FM��Bـ��/.=�JOV��.Q/���[�3F.�m�R�a&����X���=aN ��#UzX�(�t��m����F"��ӟ>�\�>�	���4�͘C��X�7Zݎ��0���1���l�lg�_#�H����\ FL�2���C5\�2�A�)�#87�*��D�L���0NL��Ҟ�Xғ�E�x4����},(׆Q���k��Frpc��v��T��j��?�xeP�jL/;7��ߒݝ;`�uNJ]Q��hГ��0e�����VCz��Ԃs|�b�y�䩬ml���;��yCj��L�`���`�B7��?�ess]����k	i�AT�0�kd���_uh�A&S똠*_���vN*M�UX�Il)��;�9��)��/�MM�*�Ϣ�R�|ͥI�� �1��Б�d&���5��HOÄ\ϩ�^���1��PPMn_�Z�Z&1�Ta}וּd
�DJ�~89�y�@13/,�вK\ ����������k�l82��5dW��  �ԎN= ̛�4ͅڍ҅
C��Hǫ���?1��9���O5�L�Wq��������k���[���$. X��BY����Ts�`4ģ�a�o�� S_�����fG��W���I�.��/=�G�~~~n���E�`Q����I��zF�jH˶����L�P��6MrG�΢ U�a1�N���.d�^)s(|�TU[����Q���F��z�	�3 ��2��ؐ��C�y[v�n�m
�\�Vkh��M������A��&U��o�\p�,L�#]�a~��@�!ƗCb�2�_�>5�+�e
���R��*=��m�W����|G�hP\�	�-�u�&-2P��P/l���Pı< =�w�s(s-1i.0����w3���P$.s��z�U4��v���^�̓�.C���V�w7!�Ti��,3��1�ͥI@�+X�5dK�~Y8��)) ^EfLs���L��`7���`��f~u�x���x��\a�z���-S�0��&�P�V;�.��*6�Ƭ����y��G���>��Z0��V�'�#������3��w�3��5h��,L}`�V[r[a	i(Q��Z;�-F.���
�o(�Ի�sH!���)T�"���w�SK���`�GZ����<��9@tC	��8S��o����䭻k����t�m�4�]�y:���]	�@N�O����U����jI�k�� �,5^��B���Q�vǚ�`�ٞB)�!t�W�29���\'���x��BKUP������L`��.�㱆�k���F6�~��ֆ�uWz3���R[�j��+�W�i��v٤�k�\��>"�[��Lspt$'�OD�d�*�����&Cϰ�+P".�D" �hѓ6,�秧���y$�_��r��{ ?y��O�ц��&��pM�-A�l��;`e0�
�dB͋����_�,n@���|+����7T�2\Vk6$��J�@.`m3OE%����`���.՜)
i\�!��"�V��b2�mQ`�`؁!��F���K��l�I�.��:��>> V# H� `����\梱�]�� l��m �W����}�h��(&�C@W��I�RfH�!�����|W�"����^H��$��L��d� lP�]�ڑ��h1\D��%ȵ�Kdr�s��q�\�1*f&��&�i/�
�E���eq.��t]�:ke^�vX�T��dkN#=+�$��Op�H�^wL�G+-�Tr�Kﳍg�¤��(��i�c���G=�'�z]���X�&�/B�}.3u\_՜��"�FE+d8�n�"�Ԫ���s�8lnn�},	gc�2O{\50I+Z�a�� X��5��@Յr<<�˽/Oe1g��|��۲��VE�h�7`��e��K�9�&>��U-2^U��Fþ�/�̇d�{kj��R���;�����w���xǆ|��o\r׮�ʭ���~>����r��پ��4�yK_[7UIi�i>��<hY���6	:�K���,±/�}~E��^*�
VQ��9/�ʜR�51���)�e�8ᚣEk��,3 � .̝��pj�:�	f�A8�f�.O���z�&�� �p&k���Q�CLzI�Tl���
�y�����l41`�~Jî�����|�k1!Z��v��Û b#�p�,�:> ]�h&��,�3�L�\#]K�Bûiar	��{8S�A�0B 5��Ηy��*�r3�6X`A~�a����4�j1����i-\FT҅Ʌt���W��)���z� �Ґ����Zi:��������l�����P��{{W�N�8�N���
��fKi����t�`�:���n�?�F����}�n�U�*`A�.O���Vk���)����E2�C���a�ѥ�#�<��4�V�
y�Z�\�U '"�a �j�9��X�W�
!,�j�n?}�@�}��ޔ���-O�SB��jzؓ��ޖӓ9=ʝ���� �M!�N3��MU���ߖ������}}[>��O�
�����y�<�� B+��]����h�SH�X� a�܄�iY�UuʰlU�!�O�����G�l�����ʠq�s��΅G��$ �{+�`ۻ�� �B��i���B.�}-,3=g�9!��<<���H��<Cy&]� ��
�|�a ����J�*�f�/(\i����ba���W��y~�SE��nJ-\��W�g���C �_����$�0Ik�
 ;��p^<��*NV̱g�T�k-����z�!��ڊ�S]���S�Yߒk�l� �A�X �c�ڨҚj^7�a�"��И�dD�Ra�e�;�S�Ui�L��9W�?}��-6�I�
%i�3_�N_$����$J~IRVW;�GJ��)R�^�!BH��.��^�(
zȋb��z�Xt�{c��WPL-�����0�3��Z��O	�}{_����o���-��3�z�+�;k��f#(�L+9\KC�z�1����L'���s�����G~,���loo �Z���ʦPOZ��@������JCyȴ�7E ���V���z�Ӳ��k�� 4�	e� w8	����œ��Xf�I?�ݭMiU\ʰ�3!A %�p�k@Fn
F�G��^���R��!��i�Ѓ�D
)0 �T��~Ӳ���ʫ0i
4:h�exs�&Ya��YQ�40W��(&�UQ�2ʞF&���n�� *j��{�<~����i�PA9�h�@7&q	..=�e�-�p.ݷ�3�����H�=;�w���k�zY��P׼P�=�����;���i���fe�<<x.�&����-�.m�$_Y���:�m�1��� c5:8���C�'?������5@z�_E�竆�e�!#��Xj am�Z�Q�B�!����T�l�m�e1��k����5Ud���<�t��}�rk�#��-k�w�� �o�&����HgsW��� �@Ώ/ ܙ+���;ՂD��-c�:{T�&�^@��*�i@��͂-�d:�$�-du}��X��g8���ṟ�=p�F�=��Y���lIg����^�
��-��_}.c�̽��R�����p��x��p�%{ͽ���E�q�v�{k�������9�8��X�?c�2(L��IA�l����R�K%ԣ�#y���<����cU������\ySn�i�J2���n]�4�
�.,'�G ���X������;������������,�_[���Gg���=�%�X���M˅��z
��,J��_���>�y/�K�����Ds{�߸-�Ǉ�L��
4�$
'*�\z�
m��h�3p��AJ������G� �"o�}V`��z0��ai3�0�𤣡Z�rc. �HY�d��x��H5D��5������lu٭A�z�ob+4La1�^G<g�<z�&^���|��gr����ܒ�х|qx$׮ �������x�f.�&C�l��vsFxFHo��ѡl�l� hxr.����4ԃ׀����g��Ă��J0�J�W����/�}�����*�I���󢬈��a>+�d9�"ˡ0�E+b��9Z@br���\�9\��'M.=��i/�)ֱ�w<��h
���d���8���@�Km �0�k�S�;��O����q��^(��C������C��u�
@8��e�y��U�n*���T,WY�=�Ek��Fa_���Z�^ER�ɲa��g=$�+�/{�8c}������Jhޤ���d/yp_�����e�M,J@���,s��\![��7�p/�}�y�Lcy��7e{�<~��K����` 2�7Ӗ5L\`��/̍G�����2O�EP�>���v�&j˗��&�B�X�Q�6�+,�G�� �կ�\V3��46�3��v���Ǚ��f_r>� ��3�CN` �����9�_�	#�L��N���F�w(l���͠G^sq�P��݉�8ʲ�h��&�=�3z����Eo�bؗi9�EY-��eޤ���)�bQ�i��A�#������FB��\�5�s]��@�y�vY�.�2��@�u-=��G��m_� HS�������4s�3NO�Z9?���эC�_wd�n�*���(��P�FWSj�zB���& ����^_+����u����U��aY��b
��ǳ�l��U C��ܕ.�[��y����B�F�ü˦�&�Nt�@v����x>�.I~���0�EY��� �Њ��ogodmècg���&�u��L�DT���C�d(!�Q�Q�w�����Š!7�#{7v�F��?���?�K������!k�>�\�(U����d<��˧ا�͵ڇW֮�a�"Y�ՐP���j"�����c��}����>,O�=�P�{��a[�/>��0�<a��r| e~�)hj%��= $u$���ߓtz,�w�0���T"it����}a4��w7���y��L�u_�|2�86*L�)�6E�_�s>8 ����6��T�~S����\��	��������h��am�A�8ș��׀U:��?{._>-&�ڋ `b�^��";V�8^�T	�AU���X��d���X�Ͷg��&,⹌�Y�#VkM�1�n������:�T@���,N��^ ��AB]5 �`%��?e�;������������x��pQl���E�{�{�i�0��4���	*�l�����v�GT��SKo��eC,��m����^��x14�W��_KX���
C�\�U� ,�9q��V/*�M�ߴ���e����'x��g����*���^g��W�`ՃR��g�r&��Zm�l�/ �a,R�G���B�u��ZkI��Üix�r �l ��+Z![��}���h�>c������[y*��� �se0O	��-��Îf%>@���}KC��ީ�h]������>��3����c�Qq��k�̴�ʜ\��&�iF�!T1E�PTa<y�ܔT�\�Z��^�e�����\{]�Y<���0�ٮ�S̗� ��e��겋��86S?�e�+��5­��"S��n���lcT�\P�yG���'�}��e���\Y�������e�s3gXb�"�?y ƺWr��j�p�L�nٖh��L�o���֖.N�8��1s@�S����e��e�oҳÜ]F�X�F�y�y���r�{^U{].��k�.yJS3JϠ��K�<�E/ ��д:I ]0L���s�=�W1Ф<а�z�+�0��k�۴��EC�Oz�� 1)�GY��b�=�ϦHI���%��`ƴ;W���q^�=��!�k�}bM�?�367��L�4���)?-;��F{c��|��H��}W>��s���l 3��Ƶ[0Lv���Xn~�-����# �k��8�Q`�>����lߒ�n��X#��y��n�MN;�MGAV8
���h^n�8���!��T��D��z5��p
 	�ށ�:Uɔ��������/l�80�m�{���N�!xzT��������n�a��O�^s�-�x�@$q<Ù������>��}�^����|Z��j�ҎW���Q:��Q����=h���-i5�����/[��j��P̩c^�|6TƩ�m����A����'Z�hEH����
�K�.����	�u³!�/VU[�P����G-_�@�����l�a�v��߶!��e8�5���/��k7U9�`�1�9�"jMӛ�Uu��d+�\{�6f{���Y���� �[Gc
��H���t��{S�jX
3�cr9�i�&<b��wJ�ْ&&Tִ"�a�z�U�Aץ�(��,�I�ۘΥ�V��Oh`k��޼E��q�L�]���
 �<��W��t<Ӿ�k��݌&Ss���9:�ظ�-E����ߕ�љ4WZx���R����T�FTN�r��H(/�|%�`=�l��a�K/���?�&�F�������L-�,3�e;���H�`�ib�/C|�CU0�.�ʜN1�����_4�k� �
Q��ho��ְe����w�F����yX[���z����k��e�JMN�ͳ)�k^$��X������dnk{cGs(b�Ik�zG�fH����<� H��S�<ƽ���jjȟ|J^�K{sKz�G���p#&�K��I���d�`^�/��SQC��c�Ĭ��w��ekAK�aD,��EJ<���ڑ_�FW*�aR��zGƽP�%ϗ�吘@Ǵ��y&N�^��a�,3ͨ��d��R�4��F���K�e/�E�)���|�?Qh�5�Ox_4 ^��L��0��s��-OsĖ�g樱 ���7j�/��o�#��ܻ��|��o 0��
���3��`Ў����� !Ә���p_= `�5��w5g��V�Y�'�J��X��h�X�m�}��9s�٦���v�ސ�m�ȿXS$4�;!'���сa17=�bZ`q�2��Ly��{ݼy`�=S�W�޴M�PM��/+�/O+�2Ey2	s��$��&��L��x�����&�(�	�z��ҁz�c�k_��I&s�̧zA���sK�sW��o�{���W�7L*��g<��`y�G�M`���{?y _Ӽ��G�JO����
M�0U���k�;�7|�Л�r,i��A� k�+�y���:�-��k�����Ҁ���#I���ȗuy��1�\6�������i��՛��9�<x��T(��vAS������| ��.T:�Ve�J����Z����Ѓ��'�O��ˏ~���p���?�ظ�Ģ�b5~�ƫ��	*��''PX��Pa_�#_zӹ��w�mi�����[��|���䝷�!׮߄���?����	�=�ꉜ�~���{;�b��*n +�f�ߒ-�6���H�7jr��y��
��_ȯ���!�j��W���ҭ`����z�I��E#_1�#��<Ua��Lrc�6�)�����d��Ż�i�fMf�"����^&��U�l�T��GB%^om�7�~���G=����jA� š������r��|B��bJd tT5tĦԮ]�Pq��;oh�_��\�*��5���Qs�B�?�x"jR���A�$IMs]F��(A1ݼ���C����m�;N$�ǲ��)�a(� �T��	�ܪ4��2�2<þ1�q��Y�r�ʞ�S� w��ʨw�MX��a#l* V�k�b���	��l����\�<kٰ�(���K�<�J�ӓ�P;A[a��)Q_PYk�g��>�bBi̹��Aك�rkJSo	s���z�=��ڱV�&�S���;�0������h��e�������ZG�-[�Ԫ5�7ל!�`k��'z�M�R�R��ǚ�u@ ����Ԫ���Bx|n��`�C������ub� +�UO���5��M�{��M\�J�������~zP�<�0��p��e��͉C�&�{�	B�e
��i�
[��&��-��;�u�M˦Ц�;R
�n}k[s���߃���0�V�-��Hsc3;�L�'���)X@�����	�	2s��p���m���;�)�=�8&�I�X�3��1�a��e���=��`N�X�<��u��#1-k�̲�т-=	q{�Zo�Xے��.�������������4!�O�6�IZ��ߖi_B�`��Q�n� �8dG�=�L֦���	=I��f��� [퇘�1��	%�cN�+�SB2MǙ�W ��c�[H,��P��@2���.�(α֛�����y6ת�J-�<z
�2i qb<�\K����2�j~v\�����G�j��P9�d[��-��4�������\h�5�vF,�`1D�̠o~�7�uqo���� ������=�O&2�� �*2/d6�e���GX�ބ��j�t�&��̷�R�A�Kg��؅4��m���G'��ܟJu�=a�� }9+��C�O��� �=��x`�n^�qg�n	n�HN!�jՆ�m]c����z�`t���ߺ�����! lC������֔f��T���&���`�7���h:y�wb�+'Ͽ�ַ��;y�^���Ĳvf���@!�@����Gk���� �ep~�ݓ��ZI�d �[̩ �e�ԫ- ( ���<���}OfgO��z�bXG��H��=z*����T�P.NNe��ְJ�g=}fb�>�1f��<�$��~��05*�B��
,K�� ��3����+Zɶ��+�x�-�.TX6�H��86�]�L;Գ��79R��k�a. �!(�]ܾ�)�W3Ia�1�Rd��P�s��b�`3^�X���
����x"a2�-X���CI �"@��vC�
����s��J�X�z�D��$u�]Mc�~�M�q�=��fG�vֵ��d04�q+m)��HCfÞT:U���s ��Yo6��,��o�]����1�������6�ŋ�(e�+�=Ǧ�.f�aN1M��Y�I	�-��b1�2� @C�{%��ee��U�z�v��;(Z�D��JaZ󮞢/%��X���`#b�e욾hyQV��~��#�D0|���fܯR��m����h"u���Π<2�_���/%��À( ^6�T2���4i�+rџH��i"s�mc�5y�ߒ��G��@�vuGΎ��2��^sҁo�ה{�jg�HT1�պ�Ћf�̵ׄi|�x�`�^8�Ŭ�O�2,��=�ea�m��D�_�^�ޚӀXiϾ���8K�MS8[h_R�!sOY������s�ΰX�p3ݳE	����Iox��c�Y���@����I��*�Ӑ�%pc:E!����󽊂_���s���_}���\�̿/�9[�p,N����hec
P�'[+s���2gо��+Ë�4�~����@<���u&��]U�����L�BC���ۊ��*�Q��\{.�5Lݮ��@�qm!�LOв���2�]��{�Ԁ:�ŏD "qar���c�� �b�6��L��vP��R;ئ8�*=�xf�wj��em��ckp�L{�eگ1(�f7�gf�9��iG�����lμ�H�LP�# 9�[���ϛ��zM���8�iN1�J�>1ҲȪ0�@w{o��i��h�9��d�e]߻�|�q�-�z�������cNO� J7���3���������TS��ί�`���ko���⡓�S�����۝�z��e�&�b֯��<� p0�d��p�H���lAl��F�}q6У��|����=M3a9t�k����>���a}rMm�}��H�Y���7yD�D��A�6��ҍҤ{����~����?x����w��cY�_��B{�-�pt�POuX��2ٻ�-_<�/�u.�����ٖǏ�����[r+���ηd4���ǟD�҅�X����� 􊬭�h���G�����P��֬J{�-�IssM6	{cEŶj�@L��E{���=PE����CĜ��m5���3eb�X��c%i��ǩ��NMC`��b�\�SIB�rShR��V.�h!�Ņ���,
#�WXc��@��kU��T�� sE�0_�����`����М������/%-bm�����&�\䩭�mzIX����iC8� �=W�AO\����*�5���3Uח3v͇0������c�������X����ԕ��C��/�ݫ��#iW=��o�����b$�f`ZG@��s��$V3�ج5UɇIh�P�2����>zdA��-�b��<��$��P�R�	#eA ���ԃ(��<j�ꅬT���Qq��R�R5�6j��2�^՜�T�[�4ܚ����zl[T�xt�-nlͷ�J:�3A M{Zx�/d���҅L.H�m�B�=_X�.����6𮖧��A�)S�a@�������G�\�[ ����Odw��e�>���03��`�A`�a>��1-a�da���9�ry��>/�[k%7����T/��#������:s�ilO�d�G�j�s���w6 �As ��F��.nc�ݒ�x�
LO$g?2�x�e?G4:�����<Kz	���9���ҋ��qe;��_S��U&8
����'��$�c��ˣ*�� YO���y�ZTVz��`�6m���g�/�4[&O3�-����4�G�Aq��XN��Y6ȴH!C��j�߿ЦߜC��h�%��pmT^�Ӳ�!�hnB��6]�M��d2�}qv0C�&/��J��� G;��s�W��r�:�﨑�j[��	Y|�04�����r?S�ckA$=ͩ��a�� D�����ϩܚ��#����k��6��dٗ�t-g�1��l�kevƼe=���T��\R<TLn9=�\�"�ՄSz��r��^��?��z�o���zz�
��AG�ޭo˓��d�Wܻ��l^3��������6A�-��)�a��	���zU����%O�>���XoKS=�w��l��5�� h�����K��2'��ݙ�8���rvq�5�5}�9����P�<��V�Yyrt$S��.�3�|P|����������o�'�š�ɓ ����x����S쪟���foGI����I�۽9�����
��f�C��ݔ���$�O&G�}�rkW��^��2͠���Ԡ\�xF#���'�뙱�U[��������M�b�م6Im����3iT
r��tA��z��U��D��l�U���o��8AV\��p��@y����pQZ'$R�9��������S��&���p�}�,Sm�D{
Y�o�=]W�U��D2�`�9ʸ�����
m��� ���&��\?K���]��{�`1��|���+�P/�&e�;b7��P�����p��
H*,���!6�w$���t�¯&Ra����4Y0��ߖ �: ��io�I\�(�J`��V�a��)���0��dsB������Bh�ӑ��3y�o��h0��K�=f��M�<f���Tװ9����ZpJ�J��Fc�x����(����p��Ǔi�\1����R�iX�VV�A�qw��rO���.C���L�^=%��e�b�k��L����	�H���A��=�4�fmC���^���8���VW�l�J@s��Sc�jط�����[��ͭ��ߗ�Bަ�Q�n�t2�ބ�
�2-�_�#;�ߔ�ù��g��n#�Ͷ%���2e澹�6�z!�O�Vte�t����>�=];�F�9w*|-�MJDa�s�Ö*��v�����`XM�[&�����9 [t���A����b������Jp6���յ��2wNO�3�*�)�G�vC5��˰^{2�C	CO����`�`�U�,�bM�D��P�XLF=Cɮ9��Q��A�����"��k�O$ߙQ�����Sx��l��ي�BŤ�h�e<����,�L�,�r�%�D�$�f�"�k�?��q�`�.S�����k
��Ϫ�A��?3�K@ȼ<=�rY#����\�Ɉ:��leT��3e�`�l�T���O�R�\id-�_v�Ѯ���젭o�G�)&dHܵ3M������{������9��F�G�2}��ӂ�
��)@�b���WV'ږK3KSG�$gK���a`G���m��k������XZrqz(w^{�3�9s���t��אO�Ϯ��-�"��zZ���&�0
#�%�ƖvҸ�E醽%7�����'� ����=�5�Ύ�c�����ƅ���(�g�!a�)���C���4z|�����l(O�<Q�Dz�� m�F�`�m�w���{r|�%d�X~�;�.�~�k�� 0ٓ�ׯ��B|�FfO������ �$m菭N' �]V_�q�ߴ7��6.�Y�_������){X��l��� ����~��ܺ*�����N8|c�F��dڗ-m�ؖ�|,�]�vHg`~��G�����g}m+�s3c�52NQ��6�֦ͦ�"��3��^ud�өP��}�U�zB3N�_\ PS!K�B���� h�\�qp���g�%l-��h:&u���9 f��;j�(�>�!s���-(�*@p6�E+�
2c�YV�.����DOV��H�ך�u��]@H���ٸ�m�r�=�����j�c��bۉ̜&�f��f�Ҏ�<=!Qд���|�wzq"�o�Z�k���{u��<��G��=�����lzgױ.�%��=���j��ː��|x_޸��H�]�B�hA��.��p����9���a�#���ԁ�H1oz(=5ear˪aVmj�\�lo���N��2�K��!Zټ09X�P�93�^��%�'&�5����h2WOrV��@P���l���1�T��B�V����PC�V�ޔ�~����a�g�~�_��	�ّ�w����4-������\3P�h�G�����Q,[�+���������i�L��*�FX�n��jX�ʃ�RC�����i=�����Pdn� S�ru�:�o,���_��+�S�!������HM4��ڐw*�Fdg�7�ʻO�֩Ro���@rJo�i!�J�g {  l�3^L���j0zNE���V���.�@��|��[���}x�v������|s�\��g�j�/�3\@�A>=h4�xF:O���<�<�k��j�c�k\_��kB��3nI?3��]6r^�m�i:F��&����bY(尭J&���FKeQ���p�͐9�\>�Q�U�iY�V��gK�.��+&�5�)�f�[ ��0�2���yn��ܔ�=7s��@zq�z�9���9��<׽��vʖD&Y�T*O��s�L�o��[%0$ s4mf6��9��M����,$���o�ŏS�8��;f>eq��zj�4֊�v��=��$�����8�b.@��Be�c���*��� a f��?ͤ�tĉG2��C.w$��4�:�	 S6�N���o��(7n�0ѣ�+_>�T�g���m��?�L�72�;�4`ccM������a�7���������ާ29���|��'�oߑ.x���S��իW��G�	�ժ�ձ0�H��)1��X�z�>��4k�|��XC��h��}S���|���`���޽��GsȨ n"}lk>0���[���Z��.t5[�A��7�����ѣ�����o�NL��>�=���#*�qp�������i?���<|�y������}�5 �����hA=s3&�BI����N��|t��fh�^��Ƥ�~� h����s�#��p�0�B��#O`��־�Y�FZ�>T]�����WS%���^�l��K��$�T�<=^��z�ha*��d>���e]���A��2���ə��m�ʍM���/(V�2Û�6�dh�(=��}��{��ҹ�<�!.d�{M��n�g�^Xz4�h*) &=-��� �!&�. �[�[&�]	�]<�'��H6;U��|[�=G���B>zp���H�ۖ��y��Ǟ� V�S| �I���s��N��7���s�!������N��O��	 ����}͡��� Ms�ʣ�hU/�W�h]zp4$��.=�z�kz��� 8���e��"�.\���΋_EC�^�������x��W5�'P *z��Rc�S\@Ya���
�����[ӳV�=?SP��}M~���r��D~SN�N��}��^����u������)������wv��?��>�n��<���O������z����s�!�V��F�5=U���U�v� �+ F�������z"׶����=��P�\�˷�����lk{���ܼazDF,��l��sR��"�b�P6*��?���4�w^�=l��1�� ��,b�:
�{���F2.�o�%����gGX���P2�" ��]����҅���{����CnK8�3�m��g�hi/<���Az	�%MQ��Il�k����.3��s6G��\S ���B˚��'�C�lPL`)v����3G ������BC��`�b�u.�4<����M`0�D�^i��,&aW�-�3E��䧸���lsz��ju�I˰.�G,&�1��P��?���w��MR�}SS�lB�.�9�N��.�O�^1���.���P��r}�2aqmM���h���ǈ��1�Y:Sc��T����C�C��T��0�N�zC�z�N�nMN�S	�0Xl�?���gj���ߖ������s9`���ބ��Tn�~M��@O���{���s�w� ����T��C�z�P��ca��>�6g��&"�?~�2)�<y������r��=]�u�Q�i�T��V�O����ʳ�S���+�}��zoY$�m����D���A���>�
�����o�?��5�aC�'�t�k�߮���h��}�u����s�zW|��bw�?��B�BнmYV.��㕫�a�@���qeg�.DL/.Z�O�=���y�����7�2�L����������E���/�G���#����9�� `�� ���ZWKi��i�s	����R٧�R�^�"M��r��"��%y͔a�Մ_F�X��ܺr��c�Xmzf��b�y�8���5 ������Tx�U�񤔹�ve�[ȣ�c�K��Yv���G���[o�<?�^�fJ=g�	�E�yg��P+�� R����ϚP�-9�P�c	\S\���sj�'t0���l�FM�N��(�YV?S��*�����VB� �?���{� K��<�9��}o��陞���;�]� �4I0X,�dڥ��r�r����KU*���eK��b  `�6����ع�v�}�會�s��$���%���53�}����{�s�����;x��_��7�:CG@'ǥLT7���r�IN�V**ѷL:V�G�BN��Ч�N��l�6[��-�Y)��57(=+h����J���q����;v�d��	��o }c'%��Ȑ�� ��>.��R�I�`u(H� ���ǣ���Z��z43�?�����~�Y�Id�ݧClp�'B>:�$�9jWtz�z��'�6�����b��6�tT�������Ɵ��_�q�p"�'{E�GV$#	x迲�>,R��:=���n�0���� ����h������JI!S�R%�i��ٕ^@p[���vc*�,-��~��!%G�ސ�OK�c:<��7vӇ�F1;�q>��#%,�~�d��Y=)%�"Y&�n4[%�0x ��X\x����K�������{p��Y�+yԛm��m5�
@�,�<w
�]%{�'(m0@Y9w���t©+I�<�XE#O���^�>I�U���/�$B^,%�&;�+��_&9�t��k��Fi= ���k��j7ͦ:q�fP}Z雔�E�`�o��X��y2���*�~;Q���X��YQi�pqM�7�jdٴ�e`��H&XΦf�8ޮ�=�����'�":<wRb�Fj�<�_�/;�'}�F��ҵ�rx��pR�5H��6T�%J��|��@#�R;�ԣ���~�Ztt"w�s��R���(���e0
�L^�;P�i�q��Z+�:m�%s�"�/�� �l��Ho��G20(�$ ٴ��Ӓa3���y�/ݜ@���ށd�hg�\�R��U�ѣGD���Jiuj�V�6t?̤R�Kͪt�H޹a�FO�۩�P	O3^��u�5R͐웃�?3�@�ѽ���<�C_�6��;y�;w��93�BQ���ą�%ℂ��s!�W.��ft���j�0��eq�]İ�sY�b���g?����9<��L�rA��)Y���ћ-k/g�M�+�j�D\�+d���`��nw��[��U�
�:���$�&ӹ�/�����t6C6:��{�3��������/p8�8��֢E�y��t08[���[.�u{���ZK�ά�o��g�\��O��Ʋ�=� �۫���#sԗ�/�z�悌���Qܿ�AR��ځ�ְ�b�N��)!!��3�t�-d�b�%�Ј��E8��=��~�8|BV�2V�]�f��Xz�N�$�"�6)����?���68�9S��;4�+:\�:�^W��t�t��_3������ �xÌ��5%%�yx�uDG,�8��t-J��p�`���_����N��]:L�ߏfۦ�;MFj>�['����µVE����B���!"a�fä�Y����$R�%�16�7����M:c� �1��3��6~�W�ag�!�rY��P��Uu8!e��1b^d�Z@�8���`2B�mRJȀ��IA[�OD�T�򜼖�>��Zw�$�N;3�l�a :���7ߧF�+��v7�^: �5�� �h�#3��,����,��Ћm���r���dH�\��P�,����C41�}qZ��{]����6�_�:�geh���?@���A�E���ްj�L���Ƥ�\���Y�'�"�.b���[2���?���]�k���elmm�6�k&8�t!�s��I����:��|�fw��oi�|l�0�Y�V�kH0c��mH�
N��ı���T�y<KS`H
J���������\�~�����<~�._B�N��ҿ+`�L`�g���O�	�{���}�C|�\thǥ,Wz�R�%����|l�0B�<� ����Y�W�qڹ�%��h{e�'�y�r�rV�u3�=�1���x}
ju�}l�\�������3mѬ�>_�c�i��� �D0�4�E�u��;©*�r��
bс�A�4�0�^�l։b��lH�Y�Vͪ	���jKO��RBh�(cZ�m0��e�m4����1*{w�ө�n�s9�񉮳L�j�PϹQ�U���$cZz��)���iV�bH�
H�6�?RQ`�{�?�4�)�T'���Z(���냜�^�A�>V�=�H֒��f�k�����1j��*I��X�L-J�" Q���Z�w�U
=rJP.��2x1�]�>F	�F��P�}�`i�*�_�A>�5�����KQ�u/�6��EL-�B��Z�@xooO�����/���������?<B�`���jo�133�%oɴ�F�ʼ2p�������������q���p�nv�fS���_�V�J��=�3B�N��h+π�=}��;<;��[�襦�k�^���&�������:4��y��ur���-2\�(�t�����^c0��dyC���HX3��z�j~�����kg�~�s��jg�;?�j��S�?��v��-�^�^9��hX{�
�%Õ�����ӡ\�3Ө�ƍ���b\�yh�wo
o��.��l5>/��Fc��z���u={���x�IX,�љ3�?�ߠ�Ϝ)�y����:�HR�{��:U�Ä�'��'���:�.�AKY셚9��h[����s�Q�&u��ZJ�� ͤ�*���ZJ��2L�T�N��eb�ஓZ���Ӱ	�]K�5	�h�HC��-��K�!67�_7��Rh9�W�|o0������D !���s�m�#%ȓ�����2D�����C[te%;c��g��K�0�E�=�J}�XK���Sd�k�Q����,��Y�!�.8\A��d���!����3��4d��Y9��v��$�16x����Nc��Y.9�m�i9v�z�4�ͪ(p"�&��-ԻͰ�2�=L�q����_�:���#��(?C��A�7�l�H��?@EC����!�{�H��h 2�=���P��'���j|�1��U6��B��F�<�`�l���N��I�#%�n�f��ʹQ��Po��	�����13�ԉ_p8�PP�]�b��Q�e��y�x�wH�A�T�#LpAVm�0�x�Õ�1��5��t���o�T����.3"�*5�{v�q����g0q#E�0Fz�$c!��^-%��&W�����T4���>��c�P��5 uk��`qs�<�ã��Q�X����u����:ڇ�`��L����tŻ����ɦ���$���L]F�oQMmx��9yO}���cF�iDbN}?f��[��,��e�_��.���0��O�Bo;Gp���;�����v��R�:h�켂��|?O��g"�}h�ۑ���I�^��ϹQ�oa��{pY8������`��K<�^T�C��	�;�&f1f�c♨U����\���5ޟK�O��xѩ9��g��%���(����ϵ�YQ��)���VG'�%+-S�21!�)6Ǧ�رV.$�hh	�{b������J�&��:�MyRf5i?�dؤ�!_R� "@�b5��e"^�} ؕ��gȄ
�������`p|BЭd�'�~*Ag2�l��?md�P*3� `�J�R�����gTV�� =�0&���T&�-f�&g0<yZ&��V:���Tz*�å42C��0Ql6cHB'�v�uh_�*3ei�v�(��٩A'��R�w;ݰx]�=����m��G�6�Z�c92���e�[YdsG8�5�_UJ��=ą�o�ʍ�X<s����@� oЍӧ&�
���Z$���n��+� P�� V�w�DJ
.�v���h�E�4��Qb/��k`=���h�dT���g0+��|��u�c�� �2[����{�}نT�Ww�U1�Z)��Ow���J�2�?�ҴHf�괱m��*p�!���)C3m��?V铚�>�Ey����d�ߢ/��>tr����\v�V�'~��^�<�L����ƶ���w����������ͧYEs�cqw����}��n��]�\_8}��Gw_��x��^�����S��_��r�|�?�E�����,���T*�_�K�.o�Q$��>��|}fP�h���**i��=�Ö�M"�p`S�yF!���&�������(�=9���t"S�3����!�=*V����ujړcR�1X�cP�X�p��A��F���2U�0&�t��&�әt��7��\>�F��j���t���W��|���[D���{� u�hZ�����;�n�-���?'�O��ǣ6��� ǆ�˗�e��/ݥ�Y���^~WN/j���-�	���WP���Ng�����|mǹ�$��
��^s�1"��4t����.�Ǩ�Q�x	S���()�2љ	�P�H)F �R��Y��1<z���0�3�>s	�{��M$N#�<���
�=���l�]gX�\½����3w�B��W�t���9��!��2dva����Ö��斗4RMŧ�)f�Q�Wq:�A���q�	 ��/�����4�;����q�d}ڭfx�&:	��`6f���۫P;*�޵h9(*ڣSS��ML��&f	��x�hC��a�#_+�T�#sp��L*��_��n	��"|�2<�D���	^�Pv�u�*-����}��yN*����~�Xjm��e��I�n��IēQ%������=Kk�r���k�T"�?����8Ta!���y`@��\ؽ������׌U_y�<.�f����A��^E�3/�)x��C�J5�=��Ԃ�qi�w�ǚ�+���.\�J��{��o�5�y*�#����tE����K��������r�E��0H-!TUyG��M��!�o:C��G�=B��>B����m�/,�[���hV���s�˵1w�,�/
k$WC�l�<�N4F4=-�^{�c�� F�֋Dj�1mA|,u�G2E A�$�$8z�������n������P2EB�c�+5�>��S�D��ޙ�ՠ�+MT�M4��L�^�F�ߋ�/N���--Y'y���N�d~�U�ҹ�@�ˠ��1	�����		�II{����$�82�@��M%�4��1|s��6d3�M,� ��>R�'QS�ϓa&�V�4[i6�_2Z�O�ɔ6����Ҿȗ�
_��t���ξ!�g�(�]������T!$�/�2�u�KbO�k������h���Y�ו�*�:��M%�b�uo���x���lb
篽�{�����S�ڶ:��n\��,m����f���R��}��X]{��ɧ�Ok�M�ԸO��h�O'��k�m���L&G{��jR��=ciڝMm�����8k�U����}�@Y���M��|��p��E|�׾�o}�Ot��\.�Z.��z���/���_�O�����E�}fvV�O��]x�>���BH�4�g/}���j�� �����P8��q:�3^�8P2u&�Ǉ6���k����L����Ɔ#��:���[}��D�������������@���↿Wm-z\���;��f���D�h���ki`�T.o��G�I��7i5�'�~�}7���u���~�˹���G�Ѹr���i��_��{h�g�c~��>3(l�ZiXw�*HI������3��qp�?�V+������-�I�X�S-J��+Uy���ǅ1�4V�
9�(���'�F~�S9%c2��q�cx$T-��2��[��/�F������<(��$|�'�_w��#�V]3�B5Rߪ�p��mA�x�؉L�Wȏ��,"�9�,�5�Ãct�t�����>��WQ�aq�Q�ur���"�	�W���.#�t^iq�8��#�k`9���M��3�WEp�:}�=LM]G��"h�!8�����{�g��J�!�J"K1��b^#Q�Y
�<����V�$FE�+�2�80�B��s�������:e|���J��Ko|g�.�ј���N.�� �܅;xW_v ��������C2Q1|���͎䎰썢Ww��|�]�{4� �kԥ'lQ����6y��*�W�=R���Ɉ"Z���Hn�aF������R���4l��m�?c�#Tw���I�un����|�-c{�A����qհ���������ͤ�Vp��/�tX��J����}x�/�򗹾.ܿ�.�x��y���Ռ�*� I�!%RK� C(o"6�ŵ+�8��#�Y�~6�_���R��d:���W?��ѓ��'����1�r�+8���_~��x�H&x�.�t�_��������*\�.��8\��nM�@��_	���@4�y.�\߆��:���	��w�m�2�i6_�c�_;�*�vE{l����0�J�ٳ 1=��_"�]B1W���'(3 �<�B��ǹS3x��i�seHo>E��� :!\��y���yȪ<k���|O{Rm�.ƽ�,$���E��Qٍ42�
n�	�'�K��uD�+�����x��._c�Ab��fU��'w�������i�vh��`��KX�v	�s ��͋J��z�:ALp����r:L$�]�V8�����	7����Ğ�e��|!8���F��g��8�Q6Rv����Ѻe2�O$��k>)%kiylp�I�_��t+g�ۥ=��:�������� �C��b��07�G����I1sl������Ȱ_o�Uu�d�̆������/��<-%p�3&�	�,͔x���+�В�����1���^#��-\Α�4 �Pa���LBc��A2qr3-�L�i9Z���>����4�;it ��]�M��zӎI�u�ǉD������~��>�B|�#s3���,:d������.3?�µKjWe����2��V�-��0sH/��^�yR�ۜ�d��O �<i�{�X9}F3�?!���n������/E����ߴK[�����_�<�޺���g+�I�6�ܡL����RW��2���+�u�����PB>=����<��k�~K dǦCBB�%�7����,����A_����F�y���&#��H�]�����xP���|�i���8Z���fu�f��v�s����g_�s��iP;X*L�N���˥��v��R�i�m8���|��{>�xF|�pP��̽+�j��$p:l�񠳐�e�f�tRG(�i�n�k;��Q��uڽ�v����a�!�m�R�Z+���x�qWȟ���������&ө������>�v���l5Q��e�vh���p#V���=�vL�'Qˈ�N_�H�!�!�j�ݻ�qUר4�Z�rj�C9�d�N�n�=�5��X6�DL�O���ZJ��NW�ΐ`$��;�o��*��M���܌|r�t�/}��%�ݎ���QEe������Ũ�T�Q#�X���/����<y������X85E�2��#�D(��������U+A�D�5Fz��@r���P:�v���P�^�! �	;?]�c�櫯С��ݳ�sh�w\[X��~v_K�҇�J�h 6t]�������D����f�Ci^�����Q� //]��k���	�	�� ^�%x��}a�<�C[�����l4�[O�`.DxrE�p�PB&��\COp��m�|��Ȏb����w�ѹ��1��Ds�:�s�h��i�høhXG"V�{��-�"SQ��.�a��~�ٍ�p��-A\|��$m}H��1n!�XB}���&��@���3 ��p8�]xBz�	��9T^J!��fq�Wa��?�	Т�����*A�5���6���V��&�M�qtp�N����`bj���Wi#숧���|>{�G�~~�he�OOԆ�����Ul?Yã�~���(���/]�IJ̛$��p��M��X��Ã�?�T<�&���z�"�v�dk�kIP��{��$�d�
���ߚ��+�$hd��M<z|}L@6�beiW�^f"S�1||�V.,cn.�Om��I3�9�m��t*���):�.���-v���<�)���,B�	��f�n��5d��E-��.��i|��S����� ���R�a��YG>Tk-��F<z��F� ���}n�"�˂�ܺuw>��ΐ��͋�����:h�E�}ϟ������𺎑�5�07M� ���3�l���]�H ��"�<X0;�b�fC�Q�sT���T}Z��iQtZ.�������<��m�y`d���$=��P4�!ӧ��tB8=����G�>:��˽m��w%�6hvR�]����?��K�x���.v:�aV����E6˦
"�����1 �� >a�0����̨�l/�e�|l�>�6�l,��$��)ҋ������$��E��d��kzRӗ'�'�C�ْM��FKy�.�AO3�7�����UU^Qz���ma��0���Ҏg�Z�沃��KP4�$��#91���i����-�ʗ�����m���/�7)����R�}A���굊��`hm��J"�����ݠג�Y!��}Q)���TZ�~���k��L;J�i�����2������c���p��~�O#���װ���S��=��R��E匔L���j҅��9����L���^���),��ZB�L�ŕ�B��+�*}Hhw�����g��r+�L^o��Kvی���ᗎ<I�Nu�P{t:g5���㟧Ǎ���|����5��.cn@pԳ9{f��彞1ψ�����Ñ�p�����V��܎�����%˨��t�~�k=a3wfZ���ak�i�8�>�������Ź���pP���߯7��:��v�H?a��c�u���F�V�k���ڛ�r�ul1K�"��ݛ���P�m��u�m�&���k��ъ�5&�7�n�y
ǻ�0�n�<#s�[��Տ�T�g��ۡA�-��������֗�Y�?��:��F}o�pd�W���G;�j�'�sǨ?������b�^4�蘮_��M��3�B��]iU�D�t��4RV�6�)�o5qx��c��Pt�]"'���P*����&Μ9��O�BY{�Rs�J���[��Aq�q�����^U<����M��a_�t�N���WE����o�5z����b/W�#I�������F���t@{;�%b�����;�׮#��ƍ;��3+8<,���:��<&x��~��W���Ïn�ʙ�x�տ�F}?{�'4�#|�՗q��;[�
�^7P�l!��^9��L��LN_'b�8ӂ2��� �`�?�̆���L���8.H_�P��lG9��k�L� *RFn*e�Ȥ=�/x%M �JB�"�Mzb���Pj�R��v?=�W���������~�C���;�{��x��	V'�>l�4܄}�?P#������(��JO����6�3�$1��~�S����0s����]ģ�x��4n�\�?��l�W�*��������{b�nP��'<q�9ܼ�F�m�4
Ir�Q���EO�}�U�C���"�ֱM����'�	��^��Y#B�=��t����K����*	f�0RGbJ:��w����*eD�w�j�-=:��b�Vv$𾻘��7P� 8�q��"�߽�����O̡7t����y�vc����I줟�����L%:�g�~���7��a�����h�j8;��A ��ҹ3(۵��Gc6��)�[8�F�,��2g���Y����\k��ￇ��30ۅ���?�r6�s�O�p�յ����ױ��Te��0��m��bWe$?�����Oov�����y}�q����\�ڱ�s#ٓ��y-cz�	�uG���,X��*�M ���c�	������:�N_�ޣ��6�r]I�%��`69�\���tQ�*�s3	C%�E���zn���<�54�geHl�쨆�'��r-�p�v�i<��⍙k��:�qD�χ�k�%a��f]e%��"���VCk�Њ�n�O�Z�� L�Y�"����Bj�S0�\/���IGq�{�#=RF.Y:��1kŘ������_�α�-T�V)�O���Z>����$vt��6 ���I砞���f"t�2h6�����"�*$�LĻ��+�y��ި��A�T����dH�)6�O8�^`^���f��l}��Hy+Ŝ�m��B�	E41Ж^\�]{2f�͓̤��ñ��6�����m]Z���Y}?�ׄf��Ӌ?�/��?�1��� j	���3�x��)^{�54�ܻ�@)ն6�5�Bgo���H1��)�0L���w��w~�����ѝO���I;��D���>}���X������!Ͽ'	���v��&��f0�8�Ɉ��~Ao�禧��^�G釦S3���LL WP������vw�*G ��Y�̓�Xi���B�.������\���Tw�?��Y�7��=|��}Ӟ`ߡE�e�M]���ٔ�r�t2{?�H���`9��>�ylU!�����S�r��꥖�=��{_c0��b��w�)��=��4
�NVr���eV*��z���3X���.ϤBoX�:����+ڤ�'��o�n�Y/|�T�9��v���X1�k�8F<�P�ֵ�^>�������b�p�Q/=vk;�;|>Q�vd�������6����CD#��f\�7���S��ץSg>8�g����^���ʼ@��Q`�����?����8궧:�씀�R~����v�|L�����-�ƨgwڳ���fn���Y|��H���4P(�[����d�D"V���+1�Z� (VU�l�OJ�T�^6zR�StAn���U$�.}%.l��JX���X��v	~���Z�t����P�X%�tB�`����!�y���}LB�ܦA��Z���9|��@���[pa��K%Ph�N_�����رt�U�LE>n"9����+!����`�9�����`=�Elr��"���{�р�=	�*7h�p�n�1������dt:���ʃu	bJt��R���>��|����λXX>�\��|g����.��i��ګY�#��)!u�ѝ-�R�P�x�t%#�����&Ѫ�$� ���}��u�XX:����m�o��sh֚�w��|�k���?�����+3KXH�'B4�6��s�C$�)F�{x�|[k븺����ڥs��so�{�˗/�������h4�����"�E����:>|�GtM�c�:LLN��kW�>�u\}������pt�X��\����Q2q%83�u���P�*.�p,J�dI���%%��@36���b��v'�cSSS3�]}FP��4ssg��֑��5�4d�\��:.�P��?��k�VR�!�c�5B�?�����S�?�B�� ����M��5�"(�O#1�BO��mQ�� ��L��{�x�W~���? �ׯ���=���'��y�#4X��w�2Ǳ2W����sh�r���Qe��m��m�9+��7�p0D@��f��I����4~M��A8���K��U@���J���q����=*�H"���y�u���57��M���2��}��u$�x�������b��9d	t��---�i��l�I��>,�i������	��(׋4�8s�Z��~S�{R��v����QoՕ���}��m���Ƿ���L�WZ)�������b�h�D�q��2�B�
3ɕ����3�@|�nt���9��1\�!"��׃��!ө����K'x�o3~� ����,�U6k���qo�����g��H�u����n��I`��m������'Z:���� �]�wE����d����l��Ȥ�p���jj���+�"b�����	c ��Š��%ŨZF�h� �2H�SǪ��Br�R�/��D�ׇ�;v"�fU�&�9���S���,i5���6�Ok��Ju#YF�0@+��X9�@s��l��]6W�?8�>�P�L�/��'w���P[ff�p��5�t*���P>=5E�0���U���u�듒�P��	��'Ot�8�9@^`�S�K��G�f�?�ݜV��?��#��3g���'6T���:�7^>�;�
fӕ������i�e ǘp������	c���K�&n40�^x�����S��ղ��m��<{�Q�<��-V>ݴ*?
�#�D]��O��tR�_�}�=�V���>��o��ŧs���L�ZYSMk����V��YS٫r�R�ʞx,�=���G�w�����gM��!�oD9{�\���6�������$os��Q�3����ID��{o�Ġ�>>� C?�cw���e�xcB�r��O�2�`�U���e�:ݪ��OwJ8H�&��7�7։#*Z�l�D��J{�������������i`�4�/8L��VY�E�mPA��K_��;�^���7��?]}��u�җw�����Aa�R	Z�7ĭ�
M&Q���~��
��(���*���sj䥗��2��c�(�lpǉ!)v������a�N��av�Pz�zح)��4Ћ�u�Q6�b����Q��L��کc���)���~��Ō:�����u���e���C8�@zsk�������e�M�N_Q*�Vs�8������y�)���]��j��<o��ǹ1�������C�y���[��'4:a�e��.?gne�Ng�������Lgt߽}�ϟ�����tf1���=̍�G�X��qm��Y��'|g:	=�J>�7c�oR�KN���ٸICPU����YF�An�UU�y��R����`nz�F,��+��g
?x�.-+�� �Z�(��p��=:��4%�ڊ���9��H���c&��[��(Q�ʗ���ڡ�� >��^~�7a���	?��"^��_���U������i��A	s����(�pp�-x�x=u�1/�v��P�Y%����	��-��1BJ�ލJ!_P{�$��/�R�����5���-J��A�#���
��Ö� #�Z�W�P�t�؊܋&,6�HUbW�W1=�c�����*̶8n�1��adO�ʄ����NXJdE::O�N����>���Q�ux?�] (m��Yŝ��;��8����2�jY�fP�Ԇ��&��(���!ڬ6K�!��̯�F�@����s$�ĕk���O��m��2�,��i�֏��	\��������34�e��c4�2�DQDd���	\��>�3O�Z��|����B��Fbg�:P#Qb מ>Ó�0P�cv.�@����4�}�W�x+��0��G���t����p�)܍��n�Ar����s��U����~8�VvW)���pee��#J��� I�2�b�@�L�2�F���OD'��m��7�Zc���}u�~:n��^��`8J�N�"Bn|�8�"[h$	O�A��%|J�._/|$�+=׹B���)����;���U�?�
��'��&T1z��kpm�1	��A�ۖ�����$x�z�AG��UU��E=�:um�+9���I�@z;J��` R�j+�+��}��g�ߩ�3N��'��'2�Z�
��0F-�����	��aU{���q��1�_T���1�~�ғU���K�̟�e�ﹰt�}�����%������N^���y��	n�򚖌U}��ǓG���7��3�+���X\��d���� IV���<�>|�]%N��Ø���T,)���\J3�c����P4���dŇ
Y���nR08�0���#��'?��Sz�'i˟={���;�!)����S�O�d����3���i�"���o.�_/�F���'S��S�Y��E�t�t��N����W��*_��z�F���� ���I��j5I�idHt�~6�M����{rO��Ft��+�!#���$i0��F�����@���H��+��ISʳ����~���8m5��;c�Y	Mc�'�J�
�p�}A�?��Q�xH��>�`<�R�J����_�$>m����!$A��������
��L؏P�=<�_��y]��K����k�pX���0�4M��*Jڎa� Q���^o�j�����D�c���w�G�鳗�?3(,��XЬm �'ӗn�S�*=K����	5J�`έd�EnzQ1	�Ì"�h�K|�.�&R��F⁠�Ly���d�g�&�j�`>i~�45R��(7k�������9<Z[EI&��U��y�:R<��?�E¹+�\��~���RJ��[t��ΝG)�ÓO����;py�A5D羀db��:һGHN-���|R-���=�Y���:y[���������|4J6G��U̮,cܰP$M�1p!W���ӬN�g�onmsM{m��̣�kO��:�@؏JMJ����^?�i�6Vה*��hJ�D��R�(?�d$�f��Y��x�[�8�;@��aLW�g����S���̸x�>�����!� z�gt=V�q��N���Ф����"�f��]�9,�������0��]�,,)�.F����Gc]�Zԋ���&i���J��01}�N����9D#��K�"�߼��ی)��f���g�V2�8�����𸹞#�d
��YJb��^�� �`o��̣�`��q����0�Jʠ-~s�x�ٱи�����6�c��@"��B�P���0⇹�}�C��q��a�ɮ�a��sQ������Ul��M�\7�mc>�Z��V%���-�e?��t��
�2Wo!5�	���4�\")�V~�z����,25���"�+�=�U;n$|�0T���W���'���(<D�5�\q�g��Y���9v^l�=%V�+/`�������<67v���k_����~�ƹ�����k)�&i(��z��[����$?O��������]C2����ɤ����@;�\o���Dr����#���`r*��(��7�wt*C�.���M�]j�JI��	��b�����ǧSVD�S�{�3(C�n-�E�����g��<�]@�����GG��P�k�L�B��5-�Z���q�����8M܏������R��^T�«g2F~����z�0�"�"�>;��������pq��h��o��j��@���t�,cu�&-��4� Fq��l��g�H[(gZȧ��݁hL�.�''�'4L�#����f�̖���H��j�5�(��hH�Ud��<)04��,�T��V�N���H�a2�
�4���*ǈ`f#	��Ye��1��	�1�� *�l�Yɂ
9Ϛ/E��!~�����/�Z��{�C���h&.�b��V	Uiˑ�|;�y<x��A�iQr���>��|����ӧO�d�\���:	%�����|�[x�׵�pmc]�C�䗯\d@"�39��J"����^�A���=k"9��3g�'����)�lb�I�9P*7��s�Am��Ih��PnM�㚑��z�Rӆ����u��!��	��u�e��9J��Q�m�y�oY'�GO�ilG)�������
 �/��j��z#CJʩ)ܜ"K)A�4��<����h��Y�lW��PM�Y¹�K������A?�eC�I�MIP��>��^��ne�r��=�O�JL1��!��85�D[&vh�[��ۢ*cE�ڟ��J��o�J�e."9S��vC2�V���k�I~_T���<�V���=��ڏϙ���2@�aQZ�.�	n%(-������z-��R��&�\������:Q��W���o}�l�g��N�ή_�����v;<8�����͛���n�Pv�l��i,ZUn�<A�4b�n�2/D��;*�.c�N�F��\<!ŵ���h���x��aJv�̈5:)���B��2�jRՌFW���|!��D�uF��r�VV�D�2�bC��D������7����a����r3	u�"�v����e�6,�� <an�_�Hd�f��l��x����4޸�#�-�D�����	@\CN���H�LN��Ǹp~�6���=L������_�5�]��J���e���Q@=VIr�U���G:iS)+�$�8y��D�OK*�����]<��J�-��w��q��U��~�N��#�fm��,��s�Oi��~y�5sG�
��|�­'������a�!9>:��N� dN��w�L$���P�Q�xt�G����«o~�\S�וw�N�V���L8�~��?��3���'�m�R��)ga&�}�����8�Pi�Um��`7[��Q��:/�K��ު�*&^W�ڄ�AF��B>{@��R�������y����o�#��
��r�G&����=�i�t��.��統��^� {؄��u�&E�ԃ�\�����'�бO�G?y��w?~�`������p���;Y4r�q6����Y��{�'�^��~����R�B���<��Q�^��_���=U�9�u�LG��<�A�3,�P��xP�k�id�<��3W3��KU� ��]UZ\8�b�� �NP��=˞R�ų����i-O���H$	�{t4NR�Y�$��`� ״QB���C-��"��8�:���68�QLЎl�U�\���b���~�v����U�7l:�Tm�-�6�2�*��=+�n�A37JEA����>�:#��f�<tb��,���FQi���^J����T�tZ�
,֟�# � (Z�5R�z�ɓ�^���(˚F���Z���/8��Bq2��Pkr���yi#������i)^ԂDID�n$�'�V �*=�L��L/d$��]-�J�XX &&��@
m�H�IyZ�d��(�������N��
leꐿ�jH�J������y���p����f��YZ�]�FQ���X�JI%��򜭴kڣ.=�!�+/��ϧ��h[����%�imm�kR�t4+gڴR�m��:��^���i97ZH08�����A�ۃ�߽�,����C��im]x�o�z�'�g
�*�:�՚[B�"ؾ�h}:u,���ܽs_�	�bF����:>!����T�891������W��'k��>b�d(�¥��%��)��w���ϟ����t����k��O~J;���6�k'U!�Z��]���;辊Ģ��{��EMXX>���],���Jʢv�)�=�����4���;m�9��?\����=�o����^�ҟ:�=�J���P�	0������*�jϘ�>V��E@%���ڴ��哲���%bl�|d,�G��@xO�"�Jh� f��o�y�ZG�\̃�V�d/��wG�����̤f2Rv������\�[�g�1�����^4؅t\���Y��$�,׹G�ܓhdFcq*�oT2�r�eHt�����  �P�6��_�_��ǩk�b�C�5��J��uLZ�z�G魫�Q@!o�g�	�h<��;�Xzb�DL�=�En5�XZH	�'��2|�cF!4¨bk3����4�!\�4��O��9�冪� ;��}��FT%{�q�C��FYR�eF�vvPdt�%��¨3r�\>��E���6D	N$�[(�k�K-�pٱ��Gj�QVs�\���˧:|S#�M��a����D؈|+�&�[�J��$����rQ�ǂ�������YC�t �����%�����o�3R�B��ț�E��ưe�?�{,��_�*�=Fr14+X{rȃ-Y2/�%����诔2B��2d���r]�*5$�>% ���kM��^o�%8t9\:}m��W���,v����m<���"�z��h�.a�pthf!E%�S�f��tZ�<S\�$ַrJx�obv��N��==a\�&�����5n�~����Gjé�y���3g��:�H���qjָ'L���IY��{��=>�%�]�����4�t䌼D����#��Mh@[�"v	���gϨ
���7�r#���N�
�lM^����l����4����iJ�{�SR`�r�>��n�{�T.��AygH�њ���p�U�Eĸ_�߻�'�� 4}u:�:?C2=2�o�����2�V&��-�Yݦ#�,J j5�0�C��=O�����,'��ϷބG��W�v�Ϲ�@ȩ|���k��1h88� (O���WPب�
\�@�{�J #0r �0B�� Zh 3��w�-p��i<���Wpe]e�e_��=���L&cvk�o�^�:�:%����qLƓ*���~[�~���u#��(��fgW��x�ഥ���q�}¬J��?h���4�=�K��&�R��Q��k&�:��\|�6�Su�%�^ıd�L���[�<�E����޸h4�U�^����'��u����l���� ��=�D���)��'���E=�\�/��E��l���D�|jA3s�RV���^5��l���5�1
��w)ʵ��dC4T�PP����Iϱ��j�Tifl:$"����kp+S� ��d4mj���053M��ןG"!�r���L�P�p��e[�ep�Uo�o���Ha�p�t�+��2���T��zEi�-i:O{_��餅݁�B$cp!���@4Ԓ� 陜��)U�Ӎ�hq�ٳ�f�[�c ����]��%���n����~kI���a������3)�����
L�D��6�W�Q��)}|2����X�d���gx�}�>^~�eUTQ���)�U	De�E��~�7��g���<�ϐ~ƫW/��`�~��5:��9֠+d�~�� ���Lj^^\�Թ�^L��p'}�:/YV������xJ�W�ӄml#H�X�UFSx��ܢ����"h�3/Z�R��s�喽7��w�`]�-��I�Q6�!)�ӳ2���*MNJI]�ۚu��k}�.��̈́��J�U��=s��i�
Qu�����6��>����\���,&�x�W��s�{k����w���!l�` ��~��|Π�����e<��k,gX���)��r>d"�?�adUy�b>(�h&�A�o3�1��,�ٝn]�B�J�K<��5ID���u#���{�3̋�o��n����t�"Oפ�qѣ8�����	>PA���ح})A��Ƽ��7��s/B�brJ�J�΢@�(���M`�Fx��6w��	:�e��˧��!%�|�� ������H#F8V#nG��U�:�����B��|�MK��z
���=�y�O�ƈ5C�0���j��1M�(�jQ�L���4�$	�f��8�ƽ�ʨ��Rg��%i���Qo���}��_f���A���ʋ�F�#St���CD}rBL<2�zH�&C�J�v"_�5�(B�����I]~���w���==�>��Ij���<�<����>��`��S�d�1٤�E �ř�����/3���JÇ7�T�g�٥��c��U�+8Z�pQi;���w��Y�����V��l���TУk?}��׏��T���D��֬���KJ���}������J\�(A6�Z"���s���O�*��w�B}�R����I�~�e�)��Ѩr�K�r��"��4.�]���M����1�& �P��/`gk�����r�e��B��7��K��Ut��cUμ�d����.�5�~CT^xNܧu�D�L��(�tH��d`S��4��T��|7���J�"Ϟ�kB�I�'�	�Q�}
���郉?##e���"�)�m®�t����4���\ѫӾ��S�B�����3m9n��!+#��3</1�M�����k�?G�VC��TC�`�S��yF=*�+����{w61�#�߫\>ĝ{�S�t�B'dr���]~^{e4K�{���$�S<�D)��ƣM������dC�_1� ��p7J�Eԕ�������jR:�}�ҝ�F��JT6��2脮<SCwX�#���6M�8�1_/�XKKI8��fͬC]�j٠��I�Y��`#[g(a�>%�62x�^d	��U��K&���%�x���լA�^Ռ�h�K�D�	ex'�P'lZ��A�:)�	Ѷ�=�	L:�� <�PJ+��R��)Y��5�C�^��+Y���p����=8����9�B�"=TR�5�^���V�O��&��d٤����1��꤅m��`F��q����H��P#H��8ȉC!��ߧ���G$8;>�����;DsZ�G�+�FW[�;�[���L�b��7���$nݹO����Lă
��w�����
:�%�g'����/��iY����i^;���,m����f�e L�(��,�tO�>��¬^c��}��ܿ����n2τ5xW�]�g����+���|�{8�	�:׭5��9�i���A���R�C���ڊ�
*�&�� X���I���2�vvwvl�:ԳG�q��Y��SWZu �ޗ��Z�p�f�<Z�ܧ�4p��$3-�����d^���2�]jK���$0r�4�L'I9[2��D: h�^C	^��NK}�P��y�m�m�ǯ8C�L�Ra�O)�s�z�]��h$�Ã]큖g$��jͣg��"+T\�)Ӌu&������#I�0ʗL��:zy���G������)�P(k�=�q�\�L*u��BQ?ߘ������9�]�h�����n���=6�$[	�s��4w����g�v�����zF��27��&��z��a���br����)W@��YI�d(�T��PPX��餧�tR�t�D,�7pG���}�\AQ��W�;�(�N�1�a�tXо4Pw�����U�<+�Q�]yh8��!&�a�������OqnڄkK~x�`���x��!�C~fW&��:0� ��&P�k��eT6��p���_���" �@����E�8D�A ������fO���u��}�3+������י�Y0��B� %$C�%��,��p�ᰭ�	�����P�Œ#d˛DP �H3�`0�Yz����׬��}_}��j@���@OttwMU��w������(�9�^����LF<X�v뫳��h��MƑ	Z}��y��]K�oڤ:h:���<p�ѯ���d|z�8�kO5�Ig�����<�1��*��) �)�}���]���c}y�A^�^t����(�o��@���"AQ4�E6�a�|���5��<(c�l �>{�3:�,�ѳ4��-fM#�'(��3P7P:��y�)���D`Fhw'����
)�>��w���x;��Bq�,-a%C0Vy�E�������0&���܍��˯7֞�P~�U�mS���fh�jYO5=���u�"xK%�瘟�⒉N6�f0
Y�������oW�FϢR[ �N�G�(���9�ʖ�dbn:��th��+,��gQ==B���M��b($�6Ѳ9����i� �*+0�++��>��ְU?�2��� �`��7���?$8���c��3��LNz�//����*ώ�T ��S:d/g��>��B/�|� 4��?4}��O��_�ދ�MfǇ'����\�U�{�3���>Ƿ��ƀs��O#(�|Qfh� @�Ҧ���jIv	�yF�:��*��z����=��h�^�$5l޲�ة�4w-�$-���28ڙ��,b��Oy.	�鷦��f��V�D���s�ly��[�O��q�໏�?�`��'  ���'ا�R�|.������ˌW��
���.�97�d��YB��n�z�؟�����&A��~g�r��*Y�L�t�뵊Ufp��:�N��g�F�������CY3����*�cU�Eg��tӃ�@�O܂�|	�c�E���dj;JX����_MQ�}i����U��=RՇ�˂��W"7�Z��cT[��Uv5/m��~���D�X����绘J9�I�H�E��J��"�Ba�U���>���cBƠ���xYA��dr�<ó8�m����[_4������=�7��C��n���x��%����}�7�5A�گ����1m@U�,�P�[���+�曵me�)ࠟ��W�l�8�?m$��f�چͽ	������*P�T̪p�x��b#\�����0I��<}��Ź���긾x�~�	DD3�a��mܷW�]��x�l�g��@�~Y'Jd��x���=����F��)~I���/E/%��)t]-J
3h�I?�J��5���Tw��h�5�1%i�R�~$�x<fjf�Z�h������W�Z"Z#����k7�r���%;?��=����������qN�>�nf��2=��"�[�܌ie���"��;��(�JH�!
+uX���#��U�n�����S��PkY�� o$��t�5i;v6�c�TÌ����7_\�~堐فy&/�Ĩ��S	�}
�<�8G�IC3���6Φ6����<HR��ҁ��I�@�g4*4#)pm� e�R���Q��	�Y>�����Ҹ����{J#IbL�=�:�:�qn:���׃ٹ �xf���HltN���6N1�h��?m�S�C��Cإk���d�ԇ�A�f�|~���
�njpϞ�����}�!�zc��V	��P!��`�s��Ҿ,���Y��Q�`qn�6�h|��I[wB�շL��L� xH�%��]9���Eku�q��b�RU.�����E�N"9�㥻���^�y�����`��;�o���[�WP;۷���_y�w���Û�%0�2p��q6����$�ް�Ǘ0��ꃇ^�˛�V��T�J/�Y�!�ŘF� 4��%|��#�RK��Ĳ$i��`�������h���t�\�	�hn|� 7f��6b,���p?3��@O����l=���W%�sOjXX�N't�O�y����璁7� K۱���և�_:�//OPb��Y4�۔N�sR�N����3~�Z;�7i��l�3�!Q��v���!���V�?@��8���Xg�8� ��ֵ<b���:�'��������:m:��g�xi�e����w~@�. 	�ɋ��vk�j	��E��_�&���*_�c��˒e��W"�y
����g����4�c���w��p�j��Kt��7WР-_��,�5t��:.�Er�� `O�N�x��:�?�]�.����� �ы�=`Uv�i&_�7%_��Ġ�<�$�g���@c�{w�d@�Z*��$�kJ<��p�#�W'��2���Vm���*~��5��SEb GL�E�Hڊv�o��@Dڥڨ��|��T�6&��h���3S��P~D3���U;,�6�x�J��q�R0��ϫ/6�e3��4�5D�3Z�����cݱ��X	<R�Ѭ��"]����,��/� ��uȬE#�S�p<15)ni�Z�����¦.EЧ�_|�LfL�T-���}-�h�0�Z����	܅U�$��8�����U��[�@�kԥ@����E�@ԕj�GxoVW�1�;��ǏP��C:q��6�oLLj4�%*�Ϟ��=����O����̓�����P�`ըӳCTM��Y�ת��k�,f��1�W!?ojJZ�+�����zV��]�_;;;X^]��z�����*���s�ë΃��إ�c4�����y��w�����p��k�>���椾�*�!΋�Ȥ��x�N�1���<����R�{�|�3���g+�E�'���ݶScR!�ז�	���_���ʚ}ƍ�W���'��E�6��,	�������l��ã6�Q
�s(����hXE�wōi�-��j�R����ĩj�oz�C�
bVe��^���=�{�13ٰ�Dc�o�󞜜�0����S,,����h]�m��G����Q���2�vT,����R�@m[B��G��U*�����>\�٘��-�k+������W��Y�`��&�<��&�H�o��yYm���<�$["�h&y��Ϧ-�;�9�ez��<���_��{�Bef�7mb)�Hs��W[�oU="���I9:g͟�8��k�\�F]��R����5�m�W�=��8Q���E���$j&MD�K�8
<�K,�T����DC�O����ȋ�=�mF	zZ6S4\b�ɻA���$�6�m]'��p���$&�n��38ρ���/J�c��:9݃ו+���J�X��V�e�b�%�7��TfVU�3����=�~���P����?�͞�F�7�U�<��$磆h�1)��椲���e3ZGyPպ��)�K�N��eᯗ0��N&�vm�s��~�7~��ٷ1j�qm��"R2��{����t&����8F�x	ϰ�_���
3�vxɡ=�Rh��3����vr�?��7������x���*�g���q��a�f�"~�D�k�.t�"w}��\s�ob����'='h%���ʈ�J����7�K�`��$�ĉE{�'bX"��h�cl�J�/���kk/��������X���`�2:�q�8�T�)���HČL��G?�~�G`T<�Dg|�⌌F}8g�<�R��y�>��ϟ����8�N����utk]�
:h`1����h���e�o"�r8�1�h��n�c&5��y��_Ǐ�{�2|�p���`[�r�F�����2�[�8�T!0�I�f#@�۳ �*��^��O���<�F���{�z��?"�#˳�k�	"�J�\���ۨ�<�w'�/�1��j�k�kQmD��w���.fϙ��u|L�����j���z�^�a�LZ��GjVr2uf�议����Y�^B�
��mmG�Kj�ͯ���li��X��۷J�|�`< ��0���#��kKr=��%���H�7�u�5t��,y��A�'t�l]��h��������ʏ�#��Z0�����	��a��5/�qS�s[E�e`sd۞"����0���8����j��%U�q<�d��`UH5����]����e ��,�=��|N]�1Z�8T�RHb���=��2� ��D�z����!NPp}s�@����y_j�<*Mq�Ō&�qq���cG��)@?b0�?z����],�\c�������p說�?r�n�qZ�-�<A5�B�r4�%-����_ƭ_@�ŭ���U��B��G��Ġ�թ�����NUMsv.��q�X4p��f�[��'����f鈟�`g�*M��%J��Y=��n�A@�52o�-��H]��r��..�6?x�����l�g�d��I>��n�ҒԱfx��`G�e��ӿձќ���Q UPm	��$�-^ȫ%)�EԛR����hӜ��5�T� ���K�tk�PI�*� ���$�����k��s�j�m�YE%XƑ�b���I�p~d����jVO�Ǫ��';.�����XF�7&���4�}	��f� ���T kjQ4�Q�&��v�a>S1]�9~��F���Ϻ�A_кE�F�>yLL��0з�������S�*��G������+�r�އ!����m�ٮ&�OOn�~�/���}@�ĈG�d�F�+Kgjڌ���d�h
T�s�贔�Ù�m��YFO��)pi\[��8}j�lsІ��d���<(���2@�7occ��z�"o��l�YUo�5��@@��Dn��<��Ï���?�gHc>�N����ݧ3l��Ac�g?}������wp�t���fr,�Ӱ܈E�*��Ï{̐�(Z|�v�Vt()?W��,�s!��"R�:����nKNr�_T�w���SO���/��[��gvww�]��ɿ�T�dc_��
�*]��t�N�����M�2�I�,��Q�l�xf(��� ��P,�g1���r:�y�)f���x���ӌU@�	t�Lƾ���e������cX� Fkm�wx(i�3��I�5y��̼U\զ�������;�>��Q�-F�6��2�)�5���/��Y��O52e���X[�bv���=�F$��;������Ē�:�
M�fF�q�������$��%"A��w�%~-�����C<��g����1k�E��aqm�9�c�nȥf�}���b�羴���۶���]���a�h����4�Ǟ��[=\e�6���~��O�N����%�f� ���v߈w�=X:/��}��n.�Rr[c-1!셌�?Ѭl>ާ0�D\n^�E4��k���������1Og8:g*Π����UV�#�"a��'�UkO����?����s�=��	��oD�RF�N�d����_��0�{VC�AT���Q�<�cQ�L���'M���� ���ɟ�f��i����t�%q&��J�ت��6#/�z�hy�i� �;��6A�H��:S� 5��pd3s�F�@"�$ȍaө���P��C&�d�$]�~�<�6���i@U.-��^9�<�ĉےN}}�# �	��9���lW\��d�tq]���η?�z�e�
���`qY>�@������5ZF�a�Qo�h���:1���m��g#&}��'�4�:t*��7��x	��6FJ�|��9m{ksT��RF��������,�n�a_��4�oC��@\gB�����Z�,pzP����w��S���Y�|Z29?G J�P�?zJ��F!�D�|A%�1���)_���K�>�KytF���#��ER:B���bk��?H@V��0%v���M���������O�>!&ڟA��N1O_y��m�fU+4�nݺe���Ξ-������ݧ>�nJ� L\��/vp��������L��Y�Ο!���L��/�'�&��j��v��5�뿱��^���(��x��b��n�6U��N��l�Z����V5�����k����i��m]������?Gx��|�a��#���&V�ҟ����3�~�C(0�,�z�*j��}�@����Sk�����ٱ��ufm�aܰ����c�xL%s�R��gV�p�0��u�Q��"���k���n��[8?.!��Y��=A�D�ڷ���Wsǉ$�ś��Ɯ-y���Y���(����η*�6Ƶ���>{��M��?);r�с�g�����̶) �^(d�S�Y��*V���!�������	��Y��i�"��7�ӣ�˵����B�&Z�K N �i�L��J�����Cd90�J-���;���GU��T��*�4�}��I���_j�Zs�cs�����d����3����}8-�b���[S��2��a�|�[����o��Z�3=(~jC�"L��ei�!��`���0�q=ڡ�!Z[�-<md���(m�j��T�V�4���Hce����/N���G��}�7��pr�����^�b��	>�o����Ӻ~7���@�/��%�1���O��[����j;P�^s*��S���k떥�j��9�J��<Kg�p�ϱq;��L��*��|�Lp~�o��@hڳe�[�0��G}P����x��'|FU�6,,��K��耘��A:�A���0PjQEA���q� ��q1:I�/3�7lH�MR�^�H�y�af^�6<éU�4��l'Pc��;j�Coڳ��=d�jUQHfm�e��f>�1�i�.^���-m'K�c�����ʩi4��t.C֬�v	���3$P����37���X��XxA0j~��@���Z!�*n��������	B�=�E�$96����]�:v����Ko}I�D��k]���X!���.t��A����c[fIE��<20��3�2H��������E|�'�I��~�������"26x^�h�9Y�16�q6]'__��A�W�V���5��g��[mޡd�b�G�R��y֨�D�YKFR���٦m+#ֵ�|^�"+�DkQE��H hK"u��E�޺}���3���ժ�{��t�`#kI�X����l�F�b"4�1��j�����46"���K���|5��\��U��ǩ�F74ݑUT	�I��rZ�>]F��ࠀ�V�fɦ��6�/ۇ1��?�6��sf�LFϨՎ�Z�'n-9�]I]�@���z�:�+⃳�#��Z��L=3��*�m�1�f}v�����O;���m'��t9\Sf�+|�\AL @��D̛b�F��u�a`f��:�"qj���س7�`�U����5��n ��_�i]�6�\#�,��4x��j�+����ݬe��L��`�Q����x�j(,��-2�:�����׸`��i��Vr�F�vw\F&\oVLvT����o`qa��:nՑͥl��|yn�fFA��*N���j��s��Q����С_�=88��Ç�:j^��=I۩��6�6y��}�>))V'��r�SM,A�t������S)37g3΍j��<�ۨ�m��+���e��<5I=��)F,/��,Nl+�0���x�3>�/��i�[6+����H��Cm�-Y����i��i��Z�4��ng�O��:34.4;��ā!��z�o�Rk3{�Z����j��4�=ݵDH�}b��Yo�.�;ϙT�6������m��X_�d�&>�>�[�g0E���*�C��i	q&���9���=�L!�@ȇ���')1�P���8�Uڌ�5k�B�R�d�H^c^^�*��u�rZ��d��aƔ��Cڎߞ���ZP�P�+A%C>�LZ�^�3��.U[��E�%��
j�bw(֊�ڭ���_(�~�c�B"լ�I��LVWs4��|���� ���9�x�0�����6�hB�6�w̉�M(�Jl]��nG3��`�sQ[D��F���b�7�&�&�����z��P��tf��E���z~�!`����qO��7�8֙]�\��套Q�{��b�c�IDԶ�uO���(sցRY�U��8�'�c������d�r��}�h`�ݮ���a�D�qfq�Gx���/�b$���"ΎO����%�3�h���P-�N���lD��e�%��L��Pu�#щe(*�"CJ�aҮ!�!���ì0����!��	F���� ����ұ���e�}��e<e�Q6CP�iT`��;�[�&j�dҐ�OYLD�D�&��`���9B����p�Q�1���[�ev��h��'&#:��[��mЅ�';���8��i�j�0�YVfZJ\�6�s���\�y}ߺh��y���Y]�'�b�FG��0����]ZK ������F�N��!�6d��N�#�_��I2GA�H�S&����23<�f���/�6_c}i{OB&\���X*��o~�z���La���ք@, "d������t*��U��#$�,��<�������1�-bt$�Do��~��S����*�ltEӇδ�$j	�l�X�?E����l�~�C��\&�H�[z��� ����r$�G�
�V}$�`'ꪮ��j�U��)�h��I��J�bɘ�IGz�kI̸G�G�8������Jz��-���L4�p5J5���}��p�Z��,f��*}H��l��D)~�̉P��q��2�qH�ȒK��1�$#��Q��,���ި,%1j�j��?��(J���k�@���I{m���~�*'����܊�c"�M��e�kmu85�gkX� �y���_�a�R%��%hТ�k�%� �C��Y[��}����;5�a>q����m�����v4���,�é��ȟNhC�՗��}��|Ӷ�[���&���qA??�ƍk�Ɵy����˰}A �����zm���R�7���,l޷��f���H��F@����W���� Kw�**G�������L�Zs��V�IN���y�](�}�o�ud�oa��x��MqVz���H\m&*Q,��ɴk�����-���d�?���G�����:�7[�R⭹3U�{�4[����L{�G����f�oq-�������1�2��L&}���`���a�@F(��8� 7�� ���f�&�����TgI"�M�\�N���R�VM݆�3?�`��A�o��g�c��`409Bgv}ae�w��1�������6��p��������s�νp���W<���C�m{�xqQ�e�p�������<_�*��k��ޝ������WƇ~nz�*.����W�B��x�]L�h�>��2I#����B9�ʌL6��j�^�ZLf�L>�6G{I�0��,�/�1���0���_�����X'���m	���@��/�m[�H��M�xVt9#�]p����|*'6/��y���iv��D}Ч�͔D
��'�o�_,��=�l2��n����~U�p��U���v�ǐ�D���4�2�8�@�\TDӉSYTV�~���U_�w"�%��p�D�Er,�4+[p�ZS���X�iQfH����5i��*���8-VU0��	�Ҙ]�>f��VE,ܚC4�@�ԃg��a&�����d��C��,�#?��Ý_�T�$��N(4y��=�	�F�>�fz�1~���iD����$Ab�AR�й�%|����1�U�*���;���?���&��^<yȬ����kx�}��b�E� c�Ci +�� ��U�oӉh���tȃ��U�T��X�7.�ޤ��b�7��;W;;������qQ����13� w�(s��Jf�H�26��l�1�Z�`��X�U?4� ��2�'�������|~��Y:߆�ް� !�V�	C##m�g�q��H[5�
cX�vق;���іB�|t>�B$�������Z�UN���̌������tΊx��ٳ�_���~0�!��*�*=G3K��9d�JX����s�{�_Ȣtq�Y��SڜU�$��_�&m5j��Ӂ��%u�M���NO���K����g��6���`\��G��?,�|z������ϟf�:���O.�5�6��M�;���S�%��u?��=^k��*��(?t��!:�L�b����.�^ĸӦ�ѽ4[e������Fq�H��%�(��6��G`,��b2��O E��N�q��%��x�1�R���l�ɀ/�3	�,AT�[�_��C��v�|���gXZ�0�̀&��P��R*�'O� y��֪�Ƥ�#�M:�n�����Y�Xe��3Zki�[[�%��s�$���h
ţS�����o�B2d��#85��s��ܖ��8t9�f�����(�<%��c6M�P�Z�#�#�s�&��F\�Tx���@��c�LUYu�n��;C�;����{���P�BK�;�����U�.����L j*-���	/�~��=YE�ImZ2^�d��_�w�Z
��Fg����c�Dt8-l�]�'o�/Nm�R�5��U�ZL�����g�AqYXE���]t�Yԋ􁗴�V�x�T�M�z�?��g���3��ct5˚�e�>@6���E�At���f�}�:a�f�ixhU�f	��\D:���M�߳x"��'<�1$��%<��~W���$��A����l�t��!nK��
����"f��q~Zq4�	&ҩ���=+l�D�<��_;\��T��y-6h1C�A&D�J�Xت����Z�Ҧ=�6�'�rFh���K��cT��'Ocmi�f�I�T�O�x^جo�b��+�K�-,b��BJ*�\��N�g��H���k�vL��VR���x�lX���ebkU�lȩ�T���h$��m;�QCkɺ�7�mUR���r$mG�mim�c����`���tӢ��KK��M�}�IF�J�pqz��X"��é��h��⸆x,l~�K0~��!�c�f�{u�&I�jt����"N�R-�ȍڿ��$C��5�=�8�������G<��'�~טt�f7�*�{��	��:�/)���s����#��>ƨ6mEK�aS��Q���.�D�8���B�6?<^3�1���M��PC�ڸ�ѸĲ-��3,�ۍ׋V�i<P]�jMLzI�G�l"BQ9�`(a�=��ǃh���Շ?��e��V����C�**��T����jCr<�ӹ$pa���,�ߞXV��L��q���#34:G:�?���
Kw�ʛ_d��G??W�;'ؚu4|}����C#	�\�3L����_��̬�����@�����_낀���;�!�G��E����鼶*5�����M��ų�k�&�L"��h�<�������4j�RP�����M&�(P�G�)H�������F'rA�����A��e��,ʗ�2��0(��j86JP1�!/̮�Y��=��%��f��=۱� �!N�
2��W�K�M�P���1����Z�c:�^߃�E�F/���%j�)K�"L�B�6�)��a&��Qm�f�T�	3�]/p��u��,fx�b#?>��c�V�w�zB�&�Ȭl��/~���mkS��HD��E�V����t�l�A�4�P�� N��i�n2���6��?h�W�f��.�F�N(�_�z\��%�.v�����o�X�A� ū!�=�8)w�?�W<C	f�7	�ߧ� �H�e�����@�t��אΊ4���t�]X��LJ��1�ݹ��9R�,V�6�}��w��;����b��#���x�
N�fKS�`�}��q v��Y�Q^�H֛2�C�6��2�;�]�����ɯ�h��0H����Q�K�hL�{r`c1�N��&z�&+�� ��BD5���ϐ���M����{�#n���<%x�M^��܅Uc�0�6����<<�Lx*�\�4�L����.���9A��g�r�TQ�x�HECHl2Y�v�D��b��s9�U@`�_>[f�+h�*&g�^aG�����}8�*�Z��4g8�^	"�M�EɴǾ�v���s��O	�O=n�x���h0�&Q��P%V�s��:w���Z���R���$��<�C#����Ե�JX�?4)7��U�% \�#��>�
�I�m���.Pu��~�.��f�>S*�כ�V�!��<ۥ�����-�&}��g��Lf"=o|�Ϟ>�Wp������o�H#�)T����ON��y�T�ƏY;x���g�D&�("�,-�\�O1��ѩ�pi-R��4@?�{O zY�_�"*�Of2�C�,��^�c3���$HP�ơl	Y��٣�3vA���Ol$F6�??�1�h8l5i��Q�B�\Iq�&��ɠ5�@a��n�n��ѧ���	Ƈ�|f��0�Q/���u�B�W���*�ji�67o����5���*��5eSY�y��(U�t�����g|��?��+��bA�;��D�#��P�ͳ�"��o���&�mWTs"i'�H�:�{��y�j�U���H��Q�ŭ:_[�X�/�[5�~|v���]���G��h�BI4��V{�g*����Ƀ}~�kL�|�A�����x̃�b��?�g6e�Za���ܡ�Z���ݹ�����C��6���t~��ngۗ�<1�Q-�ݺ�ɘzf�˫iK4T��&���8>����GE�3��I��~g!e�MӨ���=T[}�o�-di���g�kw���Q��c2p�MP�ٓ�Fǂ�@P.���Ҡ�˫�S9��,�u�W�-A��!�n}�=��RO&ހ���T�_����9	Nk�!�������!Z�Og�C���Rf��3��Ʈ+Y(��0�l6@�m���a��ĉ��NQ<<1*�s	fJ4
������k�	";�K�y`7��f6�����C��1:emcJ�k2rY�C�*ND�<Զ��ЉZ���A񲎬?a��o��f=�$��ߢ�M`�F����o��V̈���D�Og�0�e�:0j_z�+�'g�(���lNdy���5o�_��*������z�ml���[�vI �1�a�_+��Xc�^��i��A�×�6�xY��o��7�<��m,�,���A}3�,.�+{3kAwx��O �a�p(����:n���7����\����N��)4���j��&�I˰į�ь_3�_������C�BA#*�܈��3$"�$a�C^;8��B>�UrS<�4R�Np����1�������?���'��)j;EHU����@����C��#$�?A6��-C�ϋx:�*���@������Ӄc,�m0�6pxZD�]B���3#����Ne��7֯O�O�o��Ol��Y���]�� ʥSt�綽6����>c�c��1j�KN�akW	��� E�}S�q�:��h���?NQ�h��Hkw5/��{�*�������Spq�Q���\������i���l�<3L �e,�ރ����2Qȡw��3%'4;h�N�c���@K�i�p(9��>&??�~Ñ�i�0��G{����:r�yD��5��|�%h�j�*?��fҀ��a_����4`Ғ�<�&ȹ��ʬ��	3��ഄd*i�Y%��L!�l�6r�㫙=��"�:�^8��|>����l[�n�qԊ�u$��M�u��G�����$���$}�Z��.�%E�;=��3IW�IҢ�y��"D0�zq���^~�Z��LD%3��
h�r�{��>�SE��P[�ZJ@���4�I�!���j0�9,�[��-���2z�^��������1	�	�C<3�=>|�;�m��Mx	
����¶�cт	�/�a}��]�{�|��?�;ｋ �<�Ja��k3�|�`������%�����mп���#������6٥`Rg��ϥ���4ۦ�hMl�e՞�)Ci�P:Ĥ'iL�έ�/�#6��U�%�T:m2ҊV�X��m^���������͂�4)�XѨ�8M����IߞyuX罫��
�!8h��FB�1.��`q��]�5��)Z�A���\���k�)2�U�Uٴ��}�_�ܺ\=&�Rt����<���1Ë�������P�5� �|vvb����Q�F�:��6��Fգ*�_�x��RI��o��L�%"(��� ϣpŰ�壞�����J�T�ъ?�K��v���-E� 3p]���-M����4>O�Q��-3w�MM�x5]:�0z<��3�y���L4��>fܭb��s�k7��X�lG���bem��O�ϬCz��u����xo��ylK�b��٭�ڔ�Ѯ��b�$�Z�?��G���L|�A��	�EZ��y��*F��.)n�r+@ ����R0�ּ���}�	̧�K��K��Ѡ�� j�R+�C��x��>qXM����\H�%nj#>Re״YD���3\��:�6o�'�l~˶�=6���H��ˋ��tH��g��s?�?���2*�c�2�<d]ۂ�i趧�T�����?q���x��C���t��Q���	�[\m^dg����)^k���l�/�#:<��u+�i{I��햪�a������
>�}��h��k_�������#�@p6mbu}� �`/���� ?z�_�܎`���x�[(�� Ŭmg�)V���b����#����M��e��Pӈ$�Rv���eD���g��[��.97�;��V�uɬ��v�Y�ć�^�NN��|g�t�n����?�yƕ��2�ϴ	�����n=�,e��9�
�f��W5ՙ|�s��D�=g�	>c?�cќ���Hҍ�^{�%4+�H!�l\ۈj��	�=:س��4�tXU�Ѱ�[_���LDU��b��Y6ǝ��#����m�.>�3��c���Z�!��1��}��h���l��;�{w_���<n���O�� �Iͩt���Q��xo�*R�Qw�����<�#�廘ļrg��Ƀ�>�)Ny�˵:~��O����x�m��.�:X`"q��1��m�&��6�-��%6�Re��l�esl��:��Ə�N��	�&Z������1��L.�+wy]皓�;z�tV��IVR�g'm�W�4�b����O�:!�s�m�$h�^����:vEJ�+؂���|g�9��`#�)��B�H�^��$׏��,��1*�\�x{��w�t��X�� ԇ����_������G̜���0vyƔ�޺�:f�JV��T��y#"���`�˳cD�|Ϝ�)>5:��frx/��6Piw��ﾋ��;�c�Gm������&��;/o!D�������3��):L��w`���2�Z�s
jOm0�k�qߐ@\ٴ]�v��%��!��;q8�x�Rd��j'�C�G�cP-r�/����zj�wy�ӹ�ظ�'��2Q����mQ
�zM�Ķݚu��Ӷ9'� ՙ<��3���y�v{���O�^�9��;8x������f򬁭�w�,��=&���Cq�S�JWZsSLt�Z�"}�O?~��[w���g�>���m,�\�7���$��O��5/����7J���6��<B0;�A{�w�EW&xq���fi26�SP����X�L���$h�4���-ʱ�c�%��d��Ȋ���4��<�˪���5ɽL,j�[��I��7Wˋ��<���U�T �o��e�d����L�p04)W�w�Ȧ��srh��������y��=����7v��|��o�F՞��ܑy��o��6� Vf��;S���4v�l���ݯ`v�IWm����>�~μ	\�J�ӣC��qܼu�b� ��\~���B֖/�Oxc�.	����� ����;�����M�UVUe�%�Ȫ�Z��<r�f���;n��s"w��8$��#U����ZwJ!�VE���ճ�wZr!�#�����%��14l�a��%B��}�����D7`���ŏ�{O��ۺ{�b�����=�E����y��ȤD���Z�1�14�lk�(����������76m��mz��9Kcna�6۩i�'IS��5��.�k%΁�������չԽsy=�F�����B��;�A���fN¼@ie����I;�7@ڶ�a<E��2�аּ�|�KXۜ�&��;�}Ue�&�g�w$.��3�{~|n�U��y�fyG>,�`�//�X]Y�Y�3�F�H��v�S5XF���pΊ/%�u�����ŗ��8%�Ӄ�2����g���Ӏܼ���}���k��
�|]g%�o,a��L)̌�Y
��(<��(Vw������c})���7�]^D�[������ �ZP"(�0�i��I&�g/�[e�<į��+��r� ����=���n��2��ylDRG���� ��T%Q:����[�������g-\g!H�W66�%`{X2e��kx�ͯ�JK�x��N/L]<a�3���P�0��˼�0���I��.:���<�@8Aco�P]-Hvv�����~�g��M�s|Z����!Af�U\W�ҡ`��Z�ΰr�=���Bg����(V��M�^[���6֘A6y�k�/�r��{�(���dH4hOy�.f�����������_��|�m|��toa�`���"Pe&KG��JF�t ���W����]^�C�G���X�~[��@(�`Ƭ�o�7��c����ğ�cl}�K6k3V������1�Ci\����Ѯm"iˢaP�m���X&b���<������D��D(��<�,3�����>��u�ӑ3��fu>���e�33h��J;���H(�,kUj%�H�V�{X^����5\�O1K#�*0Q�Y�T:�q�;�$liY�Z����{?�|��wqv����s�#��P�>��޴J�3i'��0���	:��<��m�aIN4>�Nolz�ڶ,�7�֘���Z�2�{ʠ�$�6� ~F���z�bvptʤ-i��? X��~��XO�d<[�`EQv�L�hσ:|:g:K�6�תtjyO��]W*"n㴴Mw���ap�A-�hsqj�Z�t��ïCKc42�:����N�r,5����sZ�wh,�OP���5�!�kkȽx���ޝ-K�%ֿ���B��u���D�Y
-��f�N�����l�Z6����������� Jc���,l"���b��jm���4��wn	����8kz�|�bv�Q99��^Fx�o�6\���["��"ʘ����_�J�Gj��/�|̘|���'7F����-=Z�;U�DJ.�U���C�����Gt�0��̰OD�J�u�cU��Ɠ'�Eӫu��ghZ����f�h&�6�fW�Fh_�<��v-��ֱ8*��}�&ώ�a;����T�=D�ע-�� l�a��t;����ۚgl�c��_�u$L�x�-���<m�+L ��ֳTYf������b<31��Ϡ���}���,1��Z�5px|����_�_x?��y/;��r�
1�V�י�oX�iaq�1_������f'*L��`�x95g�?�u�,��F��G� ��M�q��w�U��Xg\�=�=hT���F��K�5hŚdf��۱�()��E��V�~]�(�gY&<|�$���c~u��{��#�Ӌ�(�Tb��v3�s������V�������C?��'1�Y��@�5�+���������F\2�m\Kƣ)�/�g�+vO:mUCÌMDL��^c��C��Q������#��s��}�'օ&c8F"=�s{��_)(����i0ڌ��a4���t��y�Y[��%�cp�`aa��p��/�� _��v��Ǐ��ۯ3�8����i`����f3Oc�SD�y�F$	"�2_��kXZ�7mBIZ
ii���#��c`�u.��qr��l����"�z�-k�ٸcmf�
���3�V���y �t6�wvn�M~�ś�`n��Q���B� �A��������6���F������3����3�Y��r6�����gU�ܸc����G������z�u�a��>���ǘ_L�^b�ұ�#ma)X�P�_m*͆�E�0~H�5�82D���}vL'#�a&��D��6V	d�t��J	��(��m.E�0����-���V�zrF�rAp�m����b�EH���w"�$�V置��Md}����6�	��(3�j33h��D�"���Ռ�h`�E�@�f��}�����Z�2�߻E �L�z�Ufĕ�!t�s�Y�e�T�*vN��-�f%�>��(
66obm�:V66�E!�H%W�1�D���/�y���
_7o��_���3)4�(F<	�>=�����@b	[w�Dvf�T�>>���T�{P>x���M�&-L%�� x�)ᵯ����׿j�����j�&�ǟ��6��!(�w�D�����h�xz���t�IB��y�HY�<;�7�m����,Z��RfQi��*7iu��c�7�������'Ǵ���"}��*��&������,S���t�����!�v';/h���8::�'޷J�7������
���1��k��<����>ϖo��%D5 ��L����&~��]�zv�ko���D��}�5���`s�6���~�R�d�� Z�,#�ʣ��{�d�m��޸w�I�	�y�8:;�\>�ā~b���o]G�����ܱ�\�zS?.�5#֕��-��i��{Uެ�<4:)����ʸ*{j6kc�?��;�k�2ð_��<#j�Jd�r6�G� ��:�,#{m{-�Z��!j�!�����eD�����=�/ϼ�g�O�p�ؽ�5�ז/��U��N||-ڕ�Z�PE,����V4�Y�k�J݀����?I����I��rQ)�5���hO	�:Uc�Yܺ��.?6�ܼ�|̇w������D�qE!���7�ۼ���]��ǫ�������۶����m�X\ܭ���nS��ThYJ��J�¢}���ON��L�nі["�g�٤Q���t��\�1��Ɣ���-�dF>Ls�U�n�d�T��׈Dmd��h�V�֖m����](಺k�Hє��G`��.>5�լ��%��a/��f��Z��>����ax�lڙ'��ʒ/*Ζn$��(����c��sm��eƎ�cwnݲ��m����5g�t��,FL���x�����o}�T>&��K&��k�\�1�r/��Y���˒9#o���VP�x�:l�G3���Kd��Ɇ5�7�X2�k�}�9�3L�H�UAh�4�³��Q��f�/��1~DN�`��xy�`�l
��<`�e�R�l,�o�c�Ơ��C~�0�r�w-��1��5�;��D �ϱp}D�<���-0�^�g�B���jj���?����X��M����+�3�Vؒw ��g��؇ꈾ#0E,C��} 8͠��F�H�*��|B^[�K�\W�Ӛە2J����RP��2�H�!Ux=�H,ˇ����@Ԕ>k�A����F�є�J&��?����Kw��+� 7{��f�x����V�ڻ��ډ=���FJ��_~�>r�v�LQ@+�I�R�lF*+y�63q�(��E籷� ��5�p^�1;����U<�Ƈ[���T|b�(��[�>A�:�:^��&�@���h�0
������L.������?�_��
�1�x��#^��A6ӢI>{��!��w�P!��1?0�}/?�O��h՚�3���yޛ1� ���,�^�a����ɗ_~��14�'`��5#˕����ҡRKYY���*>������<Dk<l4Z�����'<=�#@�Nǃ̤�p��&�O<b�H�89@� t����������}���F�0f���>�mDf�pf��tF���3��A��+���x>}RƯ��E�I��G/g2�"���l��0Z"��A��I�q��~���1���K���}<}�)�a�
�Mc[f���s�\��Q	�~��Ï�҉mʮV�%��/�L��W�S����o�ß������g��g�l���׾���5|��8�=E��ז�{�����Ӷ�MP�&�\�x?�������y�%��(���_���%���N�[psk��ݧ����~�	�!��?��v�Qk�`�3l�o�Y0p���<�l.�[��	��.���3},7��]�f�x�bX����#?�=�Gyt]>#���}��b�?'|���/S��%J�޻f�z���^���������E��va~��wwl�363���%�飾�����pk5�LZm�$�֯�4�\y�]��<������$Aa�(�b!����|��s����� s#���/��߅�p��VT"3��I`ن;�F2�Awm/>�]�[j�L���2>�~�?������\�~?|���߿�v� w�p}:�R]�)����Y���ѹxm�^\hj��'�%�2UM������Sil�K���ܶ��3-bGiĩ���4�'�����ZU��|�(bT%�����R����J!�tu&׃�%me��5ưc��]�����L��x�H��h�������D����G�{�<:O���k�����&mOU���zr���xO}Ԛn)m|B������YI�1腘����W��dE�v1����t��EZ�sW��7�9p�jQ��	��a?ڽ����ZM�sN]V�卪�i:��օ�N,]�ٛ���F�Z�FH��b��i�3t�����5mT��F�%C�}z�L��m��4���I�]\J+>�j��j�nvSnԐ.�؂Ġ2��6�Z�WOH������}ސ���қ��~̯��S���3������Xlڼ��_@nn�>m�x��E�����k���{\߼��_�>����t�Z%-4$1O��?�:x��k��>݃��P]�?�Ns���M>�r����5�MYk�x����1��\�?�yDhN��D2�����@[ˌۉ�D�F���t�}u�V�m�ĥZm�k��8=֒�sG�b܏�=���"��y�� ���lJ	[�>?hr�b
	��L�oڼ} ��8�Z{H0������� ��6h�Ǽ�a �k7��a�]�ےH5�E��@��F��;�Gr���,���������w1�vê�3�u��t��H�f�dw���-, �\"� ��3��� rc�1ʘ�'&]麂qP%g:���~o�!Pd������_�R�uMI�Dwm�M��h��� �TW��@<���&��h0�n�8��5{�Τ����#��Ј�'���n��M���A��B6aU"QUx#�5��j�61l֍�J�Y��3f}:_(�&_E�L4\/}o�G:O�xƃ��;t2��ʭM���Ъ�		�v�O琟ev{Q��>�o���bD�{F'���L���w�k����8~��;���8+�1�2�ά";�2�1���ʫ���pk�F�Nv�����l�ШJ"N���,����*�O�|Ϻ���W�3o33N� N-a�@C1�ˡ�J�UuP3�R�4�Ssr"G�&�1r�P��M�=���(B�g���O�2��ƀ�9���f��X،1�����	�S�\��Q��O/��g����&�'#�me�|��<.�a��棘E���<&�r�[���V��XW���8޴UG����	�=/
��e]k�"T�N�N2���O���fs�����y{�I��J���edd�7�mWU����?����!J���@@��>�A� A/� @����].�Y�K;�8��iW]U]�*��Ȍ�0�GdD�ܛ�z��4�LU����s���sR5��	��̜��X�`w��[�.C9�� &גr�;$P��Yc���)�8�ɦ0�ӫ��{��07G2��݃hb�i���r[�eЫa��'zb�s��_��(]E|b��R:�,�g��j�ZT-�H���1����;����u�iWD����q�Z7��naP�b6*�v=A�!9��p{ 1y�����F�4	�xku���46*��:�.6�\�LN&�@w����"Wmf-�  ��IDAT	�޼�:��9�e$��������Y�v���g*��B����8�n�#6��,��΃��G�x��)l����6R	 ���5���-�Ry\�����G$(&n��v'�c�9`��F�%a���\�-����F�&��\J�6V��0�D� �����٫��{?! ?A�ϻ�q��\ab�����OjemztN�v�N��t�	��}�E.�W�A����HC��|���'x��rۨ'����}��V��=����a�R��	�i�SԡX��Nm��zz.{���<�zQ:���M~��h ׯ�0�� �كA�L�)&q�l����{���Hß\��#H /jv�[��W�*�1�H�?z���/��QN�K���{OON6�#r��,s}cr$��|��t��Õ�^�Z��FCjMCd���CBNQl.%�R��䠀�~�5����c,��I�Xb
F]�5�SH�Ӯ��`%�Pr:'צ�f��z�q��b>�N����.�������q����<Gpv��v��g!�cq�)�8x��g����㯗�O�nr�j�~��5���p��-�u�̩�e���ɵ�>��j����S���ƙ���w%�=sG��EI��Mb�(��s�HdZXP`~a�.Ag-����4!&�;n���,���!���9x�A�B9 ����SCƟn^����O��������\��V��+��"�2"�[�8�I^{Y��� i�:��0~zO�IĩU�EO\Ś�j����S4F-CU*�$�>j�'���vQ�0uT�[J�F��%h�L� ׄl�\�������,���6���c�}RV��vC$��� -Ƙ�e|�U�F���P�������_��J�H�kx��5���d�-��)���ē��{n�0�QC%h`V�'�/��
�!�ʓϱ��~�V�T�`�k���6i��z*$NER���b�
��UAa�b���Z�m��N��<���Νh��LX_@�T
�"{�_�@�V�7��o蕘�$�I&�"�]�J��D(��x܇�gć�~��f��a� �̏�x��IV6lL�:N].6;ZRd𓍷T*��	�*em��6&H&������ƩY���/1p��}w�˵�*f�#�S�/W5aָ)��֗�bnj�L��k�I&0$��\[��F
�^G[�[��#\\d{�.'�=����21�媉�?��!���XQ*���x���P37��ZȦ8F���B������6�H�� ���E��t钞�Ɇ���z">Շ*H�;������j��`us=���L	���Gx�l�}�:�<-��\���
�����m
��`����������N�w�q�̘n^Q^7�7xj�캊��g���Ǔ�y\��D� �3o}g��M��w���_���E-�6�vw�q[@����:�[����ȶ��ƫ/�Y���� 1Cz�.^��]vv�'P��xu��rss�w�t�s�� ��4���G9�����<#x�q��T{�������%���E�bl<�ҁ�GUn� ��Qe�D�����N��W-��ǅ�jf5���k�v�D:��&�ZO&��r�+�C����%Ѥ2�e��Z�-W������T3O� �n�^B��G��Lx�h0�T��"�5iL����>D��^�v6�W�\�8_���~��赒��z�Fug�� �Y�I�ǵ��͝:I��~�|#��ʉbȉR�DB�F�T�&�����L��,��5~���VU ��g�<1�Q�<'�GH��Ȗ��r�I�1AXV�[���*k[N`�8��Y�{f����
mK��r��"��҉�t�[y�똞��ajssȲX}���|�Kx����bbdG�*��.�&U��buh�+]�v�O@���WBX,�S���W$�DHZ|��qC��	xDWt41�ث>���Hp��hW�X��F�-�4�Nԭ R�i$�*�Ϥ�S=�y�**X�+P��Ǐ�q�ʋ�D�?���m��z�a)@Y�6U
EN��y�>J���t���A� ɵx9K��$��nM���v��Gcx��:O�(w\x��	��:&�Q��:<��d�����k�UNN-N��~�w4q�'.]�I@6� p�k�ٓ��������&���C�ў �ts�KsZ���^<�����5/��"e�؉���|[�f�ll���B	l�h�����L��?�֫
V�Ft<9ý�1hp��9���}y��.b�������^��ɤ^���=�C/���S3���Ǹu�e���X�	}�c��0��t^�����B<e�^J��w��K״���Ï�����Ӏ��e��!�bI��U�F5�A��,���b!��{<�M�æ���ZU�v<1����x��ę3g��٢����֦�+�.s/fadN�N>D��_{V�K���\	J8^r8Ь���V�x��c�ھ�\y�Cz�e	�S 7T�g���5����=���u�W���t����3��iϽѠ��B���#m~��'�:���I�"L$l"�o�C�u��g��:@�$��el���������ͥ�3�D�BN�ŖN9����1gȁ���������>l&΁|�A\�L^b�z�_��-��R6����fjht�`�1٣�6�m��"�oE��r�ִ�����%X夅zGNL�e֩�hr�-n)b�+\��w�t:'8=��5��^�(]O` �I���a ��1��z���i�3H����7Q�NX�����>��}����
��\�y�z}be0�87��T��K�	D�d{풞��`�' рJ�I�*�=�b��vH�ܠR�h���z\*U��5A�cb܆�g�����jf�%#�FUl�A 6u�*�\`'|�d���F7����6 �����imEg�ã=Fl�3rg�מma���z�'{03W�G��ޗ�G~�+��d�a���͗/���&��6d�x���M5�1�1��kݐ��˕�tK�ʈY;��^��f��9��$4I^�h�5�x�ϯ��nSn�B�sA�����	RD�w���U単�[�X�$�{�gKs�:auE0�p�7XZ^W��N�9�S^WȖw�_N��!;�W����<1��W ����Oq}Y	 r��d��Kp������28(���-���.���z����&�Ghl��0;��^K��$ܸ.�����E�r�.�XR)�v���WOͽt�%�v��
����ݴ9~~���x4A[�g��:A�;��&���ED'�ags��	*���fΌ#2bЮb��BK��;8��ᮜZT�a�f;[i�wEA��a�=�E�i����7�V$A����|*_����f&�Aߊ����.rq�F�����k���Q�7�njf"���E<��C�%&�|����d�N�������Y$�9&~�pG@쨞L8������'���s��#Ip.Mu~��v�Rԓ��z� �a\ҙ�鑹G�B"����K�!d�����#5����=�:5GjR��t���(X��'��zH@�RV���Uťt\�Qk� 7���CU&PcĮI��q1��f��ϯ��ġ��-&n?��!Rey/^;��tF&�@��fCk��6K�UwU�B,�a,�i=�>�78�]&���,N8���*G�sØdKN�ƞ^�ɭG�{��׉*�~���`7�2}&m�k�` A ,���$�|���DD�� �ReLzD�3�"����b��6����,�V[�]%�t{]Ɖ r���SKm���&�\��H2F����O��L*��g��5��3I0- /�BpB�j�À��qln�3��HT�>�/�?[�m�kϔ����~�&�g���oCJ�?��yD]F�����%.3���0d���;��z)rL��V��u�q�V�"S�'���~喍��n�z	�㓌�y����G���SB�v+��8���r�?�	vOe���XO�%���/~�}��m a�k�o87b%�G~@���{T"%$��Rn �ҝ�F��owӁN�%���f��	�$=.�E�4��S�4�S�z�J���4yZ�(0]����r�Ik��9��1LH$�F���
A�|W)G0�ib�;�/|�M��-|���g�����꯹��|% >�
fDh[>w��hǫȄ���0����]�رN���ٚs)��r�Z����[��)D�����f}%6Y��C���*ˣ7]FY�"�F
.�sܣZc)W�$�N4�0[	s���
�;�a�I}�\��މ���v��t��X�xr�p~Q��.t��&���!�8UU��2�V�����ݯ��� 
(��BF�cTD��j�&�AO�y�+�Z�{��#7:݆Q���\t�͎���w�V�I�Flf;��4�hs�躶�P�$����
M�PN��8r�uZh��Vl#��-Ǯ�ځ,�synй3g���\@�x�u{����J�O���5D=]��f�i8�N��I>�ؙ5	 mr\m�h-�x&�>���n��$��>8" ��2�9�<r�0?wg^Ï�.6��\��!�B��a2���݃���*fϽ��� 6��g<}t&nh9�����O2��,���h��Ǉp{ ��8� ���Q5�:ݺ�}u	63��z��x��VƜ�?Vh�7���5��m��Ֆ�N�v��lE�K<�:G�3�ʉ�n�6��#�b��p�\�7���0���6�2F]'*_���3��0��t_��;��d��\�8#b�W��S���S�x�>���9��{�������iG��A�YC��^���_���ݫ�r��^�c4!��]�*���v
ӗ��Ig�D���E&a��w�b�%bh2�֚��$��A�F�*�Q9��_@�|�,�\��p�@ts���i��$�A��N]���pt���X�~�M�U�����Q�(�q����L�$#/\{���	��ƚ6Mό�6p}�5��}� ]�')+8Q]�q��|
q���ѳ��~���XBv�z�� �+��8�{�����~��}��+^�^�S�R?( ����VSL(Tn��Yw(���G��/�����0αm�G������T�i����z|d��+�^��;�)�E��F�@`t0$�:�����v$����6AX��!�n'F�68Ƚ��P�s�T19FR��a&��Ϟ���k�p�����{{�r�����8��{�'	�cPk,�%��mrNln�R�'eHR~�;�b�q���C4�W���Z/&���JY�O{�&q�9@g�`�풝������8ZD|�I�ĶS�D�jG ���j���?����؉Ο�4�8��r�l�$F��j1Vɞ 8�9� ������S��Q,"ˌ{v��V6>k��P�Wq��S���8�B���zL���ȕ�@Bk��z-!��W;�.�v�s$w9��9r�i艳��a�8qR�V���,"�k��X�Ȩ��I����B�i�M'���#�!��9�*�ӆ-�0WEx���gJp���	f�'��_�\�aj�k΍�?z�/�q7�
 @r�4��w	�1#�`;w�`čs�Čz���H��T^4"	�%V���]��=C��;��6J�ȿ����d4�]��f�.�� =���d�H�o���X����@���:����F�)6{�%թl�*���Y��Qd��tJ�~d�˵©��4dr��[0������=FC�n��� �W����q�45C��Zf��%�SZj�����at4��
�,���#6�2wڜ(��MN��b�c��w�>^{�3zb���	�</�C��VE����1��q��Py��I��X�Y8��zKO���YdVD��l<�V��Y9�:}9�i�ze~�����(i\�k����vT�C0�h��p��nO�_�a�P�����TG�[�0�DsQ����Th�j=^���K�ē�CPg�n������� �v	����J�n�\u����D�W�-����v�H8E��A�O�"�$��Z��@T6�p?D~�M�bH������il�v���b&5�.�X��Z���R�/RC��]����X`�+�B�E����kH��adrw�dPh<���~V.�L6���	�6���y���9�bl�> �$g� Ɓ)�L)Ái#9�c�G�	#������!�g-&��Z��qy	d��.G��I�	:�O2J���`y{5&�}�fUm4윘Ͽ���n�V!����Q$"Q�E8�b�6���E\8���إ���#6M]�%@1{��Gð�&�uU-p����ea��$!�ˀ)�&��"�y�>�����o~�w�.w+K�?wQ�H��->���"��Η8���?�3$���O*G�r8����1�H�DBa���
@(LV�WW���U�A����>��o`:Ľ��G�f���n�xC�
:�,�2g�T�� �&��U#��y�/������%�Te�Օc���q����GPl�� iA��!&ţM���jb+q!����� �v��x��Y&.�j�`?����ʪln�b� Ip�mf��̕���y�2�5���k`��xcq4�-�tJ��8H�^X��[o�'?���69�|�j�̲	K�I�lœ�kdd5LO&Pe�ٜ��M|�뿭@4�_D�E����I#m\D)[G6WQU�G�n�;�>���ǰ0�|eB7{)��$������.DV[4�W��� TΖ5�U����~$���~Ģ&�k�Z����u���DA2�u�5�Ծ�`�v�K�=籹� ~��F���׎�ވ���\�xE��<|� ����q�(ǣH0!� ��u�BUO��V�3�!>ĵ�@���G� �C����@O��.�mhọ�K������q��65��xaO�7	��;\+]���3&>[0(�!�Sc@��z�ۈG�NC~&��1������Ԇvw���|J -&�e�	�~����8���E�slkG�jw���qgm�@�s�up��c4�S�:?�6��484D,�{Rn+@���4S��I�\w�t�^��כ]���a�7�9A��7`�\D��Eˬ����X��sX��$�=��t�����0c��[������q��� ����i��`v���B��ʕ�$�V&���'�m���O���?��Hd�I��:	� J�d�˵���E��g��aH!�+�c��NI��.]�Hp{���g�B������&����/71�!�EP�F�|� �F���<	r�x����&Iʙ�s��*��� 	�IKo���Rj$Onv��z�ASu	MZ�u��>�J�FE�j�.�ۢs���ηq�x����;�Q+���y��1�G�D�O�i!!%�l����>�$�� r�2��/�����93��==��j�J�Y��D�Y�d<喦�������줓��qu����N4��$�(�s�(��(���.������C�LD��ص���4U�[<�}>����Ů��y$1��f���	B��I7�������=f���d7��s|lB����ν�
��k���c(b���9�y7�n4�'��6�E4Q�$��������K9����#N���SG�!��RB$��(�H���NGeh��mu�����H^P�yY�&#	S5M0H�1��!��~,���$d�jw+7CbC����w�/�����$q�-�=��:�F1���GwkZ�(��$%�����PN���v���̳E|��"��[��.��c��|�q��bw�}|��_�xU�JU17s�ѳ����,d�1��nsJ����N� �#��f�?��چz:�j��#�_(�t���@rb����?Tcp�͉J�ą:@0b���H�?-�� �c��]��al���T���LR���	
V���j�p����Y��U���k�.��J���)?�c4\��a�,�h?QS�2�g 4B���"�sw��-d���3y&�8���
�d)����\�>d�e�R�����J��V�3W�
�\~�S�1D	�6�����>�\?ڴ����%�~�r�S	���������@���� ��/�Ǖ+��Đ-q� ;�j�1���,��
�D��_~=8�,�Z)�L�F�H��8Yҕ&'�b4.����(���N�Jf8����ZP-r9Aw�`ҋ;wayy�����ֈ���rBʍY�aj���SS.��e`�	:����h؃��&�<<�b �&X(���p��u�fV��f}��kpƣ�q�!�\/��
U
�h��Uk-
G],�.�=��U1�jg��,u�2pcW&l�g	�w%��L*ŠB�	\N�$؅��?S����
���{&>���&7]��uM��g��zR]-��|$���=��dǵ�s��&�����+�/;Z'�bR�{���H��m���F�Iq��@�;�+�.=BQ���:r�j�LH��T'�"Ǹn�C4G
4�m�����[`��cn<���I��#�a����z�!��w�<ǹ�q�F�t��h.\�MS���{��5pz��DVpȤn�M��!02�Z�S��<2���>��!L�"h��kFL�]h�;�ۢ��A���1?ND�KN��E��m�	\��SM�i����U����X�� ���R�g07����Ww��Ԥ16��b���tURDN�Z$iJ�H�����/����f`���0��Wf��@���֫7��\\Ο' �0��|ܧ���>=4�Ia����g�I�J��N��Ht��VM�F��|��?NPoCb6��ERK��������$��U#cMvW�"��e�E�ԋpd���1�dr����l��{!2��'ҩ-����{��&�i�$=�穛8i`{�C�1�$P�&��bIkԭ��rJ#�rzX�Z2[p9H�C	<#�9;�^�	����Q*6	j�sc�qe�Di�~�.�An���aor'�Ž����씇��`r�r/�(��c.��Ƌx�xg�pa�����1�$"a�I���O
����8���&��α�7��|L�VU h��Vzx��`4q��ǅ?�����ŇqM��SD��ӫ1�����k=�2�hr��7�ZK=>yF�5�V)�#��ٵ!6z�kk��!���g=>��F�J�N g׎�i�i�Ӗ�؋v!<|�VˋO����X_Ւ�[/����8RGi�S���e�X�����H~�NF�!a#8 YK���pG<�MZ ����R#�4?�kC$e}��ե�Z�V�*Fb	gr�N������|=9;F���c���Ġ��1q��|��D����7q=��^����EП�<%�w�mi��*�|��9��m`S󚅀���j�]��R�dy}^�A����I��q
��VrRR��vSC5B��o���G�ŉ��&�ϫb���q���D�k�X�C��T����5�ZI��}���S��^���[\Gr��8��D�6������F6s���;�u�5d�$�W�%{ku��2l��Q���>.2�pM[{�H�\1�ۀ�����H|x�3������Mr�-%0�O��ڬ&7�ҋ�Ӣ�_O�1'�r"E�'��n���e�@|����@0�8YJg��z�q1ʵ�&����cZ�^/2!����e��Fճ��E��j3i����%2���t*�j��#�2����Ȋ_ܹ�#N�̥KLE=^�8���:-9?�F*��3�U��0t)
WK�񡵯>���~��t2�����bR�� Y&����vX�TT�V���{[��9�k�*���kQp%v��f摯vp���ep�c$>�'����c5���������y�u-#��ј�'I͠X�I������;�[��݋���p�޽�O,T��\%ls���G�B>���sl�'&�*�9^�� ����q��?�s����?��������I��^{�$�4�=�֎AY(�"0yˏWd����'�ĸ�f]6&���w�2�$3��P�װ0c�`{�)f�~�˻���Ň ��ΡC���BE<Nl,�ݔ���i$�ZFbr��b�3X��`�ar!Z�{��e��|�lC哒�I�;��շ^E�k���C2� Z�"&�������uT�3q��y��	R�Y�������p��^���}U���|]�|�E�1i=�!	^	��	��U<#�}�����R)�xr��PkE|���k���*�a;ff"(���'���߄�Gj�	���DKDg+�}�e@i�����P;.��2�z�|g�6!�Bb����hU�m6�e�R�������MI���m1��Έ���vx�s�Т��`CkԞ.��Ɗn��Z���dU?���Utpn�@�`��\���� h!h�:H,c�IC��4�4{�����������P���Ͻ�b,�­��xv��{\?+������	�$��RV�*�\��Y*r�����H��1��2�t�A"{x@ K�])�W�t;��,�F�D�c�"v�_�գ:uR
/�N:��*J��u�ڪ'�������Zllb
p���>�V�1#��&縄�\c��Z��d�94�4�����v����Nq�J����8�r��s _��"��ʄ��[�0ີa�i�_��So��[I���]i�ޓ="��no@*���[���$!5��P�F�@� ����}�)u���-�����[1�y68(<ǵ��$��w	�l������*��M ����Ƌ����f��7o`h�cv>Ap�ŽP÷��
��^��	���� <:"�2%��pm���J-��9��y��
�{����%~Nۉ{�����e�:<N!�0g�a�\8��{Im�]{+�+\s{��?���H3��ʢָJ=t-_�Xrg��L�Pm�ۯ�5R�&2Sn�5�^�Zl��#HM���i�Dڬ��(vw601����%�a?�ŕ����������bq���K�dP����E�;'&	ԋ���
 12/J����HW�����I'Q����0��'O5^�rA�̵#����7E+� .w���~�r����O��mL�ܥ>R��c$�Ҩ#��f�8�8T!C ��:cȥ+8:�Q?hQƐzC�r����q:J��bP-��F���2����8���z��aJ��{[Jb�1��&�e�$ˉ��*�}���'Op�r�~�kń���#0��I��lS�,E~���� �#��q�b�96��g z�ԪJ}���-���<�ݹ��ҷ�.ސŽnk٣�+��r6�b���e��a,k�q��%t�),3هܷ�M�q�n?E>���E��W�c����یW=b�&��Im� ����S]Q�f������O�I_�ɯ��֮�`'
>@��$C�'�I1)#�-�6�g��"sq���I��Z%��W��f+��vA�G�Ec�X��o��M�`�C�DDzC��ۨը�� j� ��O#S(a{7+F�� u�	1�P,��ػR>���`s�9bDk	ϐ	9��Vn��}���dȘc�	��y��f��ځ�2�zfCQ~�`L@�� �[]}n1��G���yD�D��9�_zU�����	%���q.��|M;e�>m{���c����?zR$+V���A7d ���S�'ג���<{�\�ꛭ�v��?b��\��lLQ���:��\�K�J2��o.i�D����+3��?�s&��|�Μ�ſ����w��9���rO?Cj��.�ݩ�=>�6V8���"J��V>��X$�k�|x%&���I�Jm�T|�LY\�˕��t A����q�q�ɨ���HX�.R�k@ԁ��I������Wq�/A��DH�˵�&S���o��t�>��kgq�0�Gt��fh�$�µ8������qs��	L���+y���a��It�\/�����qѷ"4��p��y=N�3�taF�T������Zi2Q���羈�9ȹ��ⵛ
TK=�V��5�:J�˦��ZWӐq)�&H�q]��(��c�� ����8cj�f����Kx�A븘�8m��#�,��淑$�e��Z{Ff�w\a��u�oT.	��c�̵K�1�|x�<f�ݺ���>a�4���7k�H�|#�i<&9�ݧ��L>5&����H&���o��us�S@���^��`Ϋ	���1�K��!��(����$��<=�Z��ً�N\"��:$��:����cU��m�8�
X0�<*�*�k��&ZkGx��?:� ����^�����z	�D�E���;!H(��(Hf���C騟��JD��)�kS �E��'ZD.5Y�"�*����x\�3����KO�7��#D!|�~����h �X��L
T���n^<�ן/bwaR��!�W&f�v�V�$��6IZ��$�zJkut���f,Q�H(ծ��.v�}7�Ӻ�N�k�cm�ԅ�!n�<r�&㘑�? CϤ>���brl��ǉIU��\�.O��O��q]����Fg�k�Xz�K����|�&s�;�E�E,��𼰍ɨ�W�nd0;3�ݽ4�	~}e��	�Qt�䦏�)�x�k��u��p���=����WP`=�������x"���Y�G�ǧ�:�d	����^�c��#�����Z�#��q��HZ�(��Rs6���O4�\��*�':��B)�9�SM�ɱR{G�Zn���I@=������|���\�U̐즏Pn��!D {�w!62���[��X�=�j��ڤ�N����$�
�l ��4q�9�K&�(q��Nm��X�OO�	��C�����|��7��R��' �u��Yoc������W�����.�ݟ���/��z�����(�}ϗ��$A���£G��JNNN-�0���N�{ۚk�Sb��X\oO8
 Mm/is_�R�?����`.).����"��h�J�����e�F��F�5�U���	��	�$�Ϟ<�\�0�3π�YB��-I�y��S��?��v����s��;��3�[Z�Q)�s?������'�	�,�6���@+��F)�.c���"�?Y���0�ĕ�
��r� ��\�T��-\��ڸ8<���֊�h�4����ME��ĺP�E\�������v�2($��	� �:�����Kp��e�1拪'����ND5M6�"�݀��PV-5p-&���\/1�H��͋.Y���8��!���Z$`�;��5`8�J6@����^�jn&��h��"̍&B6u�`��_O�O�E~� C��!�y�,�V�2�l�	:���M)	f�c"�[��I2�o���bz�g���(��t����w�I�t���	a�j�~���j��fГ�������/&,�;;����c��g	�#�gb�����b��x\ G;{�+�m6�\��%��2척B*�,��hv�-Zof`����D�+1:Š��SU��[���a,�఼���Am����T�g�^�{��'\�W�_Ƶ�����M2�k�l�] p31��06�C��%�Ki�F`���!��Җ�r�3��l��a�&#�;�7?����:Ϋ0m��[t��gWNo�?�_�3h���q�5�w����u�z��Ylloo�'
��t1�䵝mXN��������9-��vx,~������/�]��Y�|.H VRP$��+���U.�&� S-���L�8�Qđ"`p�TH�p�{��I	uq��W���	*�>�\x�}��Ӯ<.���c&1��~�����h��y�_�����:�'�i�������@AB6,�1AVl�<�V�O؍W.����[*�`w1��0��;���_�N�݋u)�H���3`�|c^�ե@:f�J&���oc��e5z�V;HL���_��V+k�Hv�2����6��u0��?�t���.b�������ο����p>�����|~�8��P��h|:���%���B�! >s�&B�s(w��7����K���z�R8�>�"�+�n6PI�6�����&g.`��8u7 x%6A��f��+A%P[����X��8�l�pB@P%��=���6#�=�11����#X�KR��?�6��苗�Xb���e�ȵQ�>6ٹσ.4-�$gP.�Lw��A�O ʤ���}+E �dT깘 ��ݮI睠��7��=g纵b����_-ƣ������H�R����k7�dG�QNL�$�L.->st$�qeh2Ƙ���fvi��nI��	�D����	a��-dv�T��c�U!�wq,��C�m�;p�g�;Z�b��K*w��H鑍q����/]��󏿇�_�B��s�wmBn�����*��Jt�@2޺G��}0�T��3L�}$"�$6|�8�-c��1��T�k[�}��̓���7�����2�]g|;$h���T��۷o�i��>i�\_��&�3g�c46v�$C@$�X���	p�����,2���n�t�5�J�&����Z�z�}�&������z��_~GK=�Di$���tY/�={���s*=��o~�:�e9ǳ�qDw��ZN��ȧr��f��j�
�	V||N�60��ŝt��s�H΄�����9���`�����q��U�-׏1==�*)�j��1�o����(=~�.<�KOa59���p�c����L����{���Z��(�z�)�Q��jQBc#>�Y˼�4��|/�Ȳ^_�|	��>q%�ȱ���>��w�L�Լ>އ'�%j�it ˱�X����6���52@�H��{�I�Qf���J)�A'ϑkpZ�v�#�{558h�~��w�|!�-rn�d�E�~���j�	�J$�G����w�j�o�{9�'��e1^;�%}�FN�s;����YI���e���'yD�ټ���h��9V$g3��u�딤�j�B<�.�c&I�Z{�4I9�E���T�(����6WbjB���m����%g$��UM&7Yc����A��o�������t@4�u�ހ�=�$�����Lt��	�d328��P5����K��;����4kx�=V��a+��X�ٹ�݁&[�n�;DSD��ۈ	�l�a�u"�#��M <Fm��U`��P�UjՖk�c���$C�d�+װ��#���5Dld>�����͚��E�z�-�f�df\�yU��|�����ȷL�Y�Z�f�זּ�njH�z��hm�Kt���z����+�E�p�D,��Ƭ���6j�_�����������L0ʄ�A;����Q�.�l��GX�0�^���W��V�w�(��]���וa:L�8���0�l�nq��zŞ˒y5Nk�^~�%|��66������?�"����H1��p7�8�"�fC��z_�#Dk��s��9��ق�=�?��M�a���%ܸ4���(�w��ɾ�D����=$�3\�8�0��#:;�/���Nu�c��N�D������M̞��7�[L�nnb�?�F��*���D�Dt8��V����*|�c��UF��ڈ��Ns�>��M��6rפzs�~΀���א����4�P�\��q�o ��X,Fxc&��k+�h�6�kV�98�\;��v
m#22�/�����>jq>c8"�?ӓZ�^oV��c18[��g��Z�	�����.����ρ����$��:Z]����=�xDk	}~��9g�Ӯ� �VG�2řBꂧg�s.b�Z���[ȉK��5���]8K`�qI��="y�^'�KW�bt�,�VqP`��2I�� ��̼I���Ʋ:Br�NE�ۜ#;��A��˯�M@X)r��9��?'L�'C r²��C�6�=gc$�D��oL'�kU=�v`K���Q�u��L,'�'FTf���l8�4 t[u6���k�f�����/��d֢�w��[C�I,p`0����w�����zuIn,�Q���h������G��?3��c{�!n\���W@��O����b|ԇc����y	2���*4,RP&��V[lԌj�%vnf�s�I�r<�$<�E�!�����10�[��kH���ך��xT���'�c��0?5���.��!n�p�{���~�%	�ym&J-��;�j�	�Ϣ�qj��4I� ��F��i@ ���!B�>Z����/�_�1�f	606yN;�#�(�_~r;y��gThYj�+f�4!͉�ϺD���g��Jj���A�3��֞�����ݎ^�����J��=!9�H#�%�R�#�uB���C�M�)h�5(5��aO�>�v+.�����\/\�I����G���39�_��{x��E�$�F<�%���+r�J���AV�3a�;H���*���z+e2���I�O��FUSPZt�$H�-(�O����v�BA�v�5�GI�H��i实D��믿��u�$��*IC@w륗��t��_�������:b̡����Q�,Wdr],�	2�z�+1X:��W��v6����u������!b#Q�l�\Wo wX����x_���~p�y��
�(���xP�����!�$�-�11y�p~�����V��c�Hf��s�Q,��Uw���̏uX�'�K���G��%GN��'F]��'	�̵*��d�7���;�Q��<
	C�q� �SJR�8^ɱi����9^	���)��T=��/Ph0Y{"�p�+pҥ���EWP��j������G@	����zju��\;jUu�``�jFА���Hm"�x�؀(���Z;�"��ol7���3T��
^^�` �����pKW$���I��	wy���ʥD�yD����Zrt/��LW�&����m�\�U�Y�˥X�uL�Z�u�w',O�aW�6A���D���n�"�����s�h���U�^|�	&��;��	Mx�r�(Qcb��	dv�111������8bn.@RŠ�$�v����c!�5x.�^W|�O��ÝL�h4ڑ�-#G�?;7���PͯR9�=m8���x�|�����J���f���<S)��K�����2n�������ɜֶ�jY�+H ��g�M���g(?���L�L���,@�'��L
.�e͗�x�$�r�026�gk��t����V�Il8Hm��@+EnA1�,qM����}�3/��L(�E!��A����!��!&Gf�L%{�[g����B��q���Vw�D���ͪ�?�&'��}��}��AdlJu�D$�%dm^2�.����ߋ��f�n@(��rS	����j�^�af~�_�|�u�����o�:j��d�[K�0�#�)�Uti�D�I DBS�l3�ڑ��b#<�8*$~S��Ϗj��3@p��rY�(�@2pa,�t��EH��{Y�	$G&8�-D 9��}���߹����}�*�p���������=���U:	b�>$2�Z�k��vOJI�ؖZL�I��_�H3p�3�{�ˉt&���]����&%�AO[_�Q�ַI���W�S(�[ʃ�z�m��Yg�C�I�����:T �d�����ˬ�ܛ���>XQQo7z��S����v�> Vr��sx��Jr��LDs�q��|N9M�,e�'���z�ΰK�`�Ճ��]$P�&�Kn��dR���܈D<���+E\�p����G5I��"c��Ň0��0T��v:�UZ���494�ky�N�`*1�1xgw��(���U&���1Μ���V�ۚP�TUI~�$��� =&u�J��DL�ND���ӆ#'�O�-�B�Rk�ObX͟	o�$����38�����Iv��[��=��*Wn����h����E jM���ź	s�s8������6�(�8/=�0��Ft$!h�FK���4L=鄗��&�W���󒇥7@r�Ǆ�	�W�y�H�Ț�����ƘXG?����l�Uҍ|��5�F��EH_|楄IDP^n�,�Mr�&��Dz�#&���O�����nv@X��)��A�:�����F�3�LNN��v21��I�zttD��̹s��
X&�	�|X83�'�cЛ������*�׮�p| L@�jk�2ѓ�s9���ѽ���HG$���v�Y��7��M� ��+�-�*�x���mL
��L�@*�V����U��wloo�x�x���_�2�z���X~��<0��E���j�=~��Ի�C`Qq�J����i�z`h�hR��~�0���<��}��;��;�z�9�¹#��̧�X"���#��|�r�����ݓ�̡xFl8&1^YyN��E4A����� fc�2����\��r�̍G�&L�G�-lgi~o�^!�H��{�Q-wIL��$p-�\Ʒ���I\�vU�T�7��GGT�;st�2G�"kD $��$�|�]�=&�c�œz���h��yB�8�p��ܞگ��~u�;��-�b7��Ʊ:LL�G*:����ٍbt�:�H�q6w�E���]Mxr|�FU@��	]�xg(:Uu��l>/����%��6�N�p����u�P���,�'3[Ы���݊h Z�0>�i"k���cz��8�##aLN��BI{��#�j	fg�uߩ>���0���o�]��Z ��뒹Y�-�ԭ6=j5#�-�%���نL����-8��%x!����ۉ��kM�/;����XdP����.�LF�)���2 X˖Qb��D�h��6[rM&��M(N
c.o��=�,/�M�G�"�>��6��l�"��m�Ts:N��2�����Ǆs�%��@��ȄrD ���p5q~����&������uT��7�k]�t����L��֠#�w�
y�)α�A��K�	�OX��ٓ+H	^�����E�?��	lrh�`���y��]xBv�I.1�J��tr�[C�~�����Z&?�G�1a�h/�*Ѣ_��N�o�l2A0�B%��}Po�ӈU��X����$��dI�ҁ�Sm��O@�K����hM덆-��p/���^c&�lJ,�8?�8�R��v�YT�o�TO�l�Z���P����I�d+ө.�\:���b�'����<��H���-�=A�e�e2ٞY����P^\�x�|B��@"���~�Whp�՘rR�k��s=��%��'��)u����Ԩ�{E:[ŗVN<�R\NĄW|v[>=��- ����>7"Kbc�v��&ـ��'�mR��2��	���'uS��[ȓ�P��d��z.	��Cf��>#�n�VG,�F�Ib4�B����v���q�����0v����	TCX���H)��$+����`"y,�V�-V#�D4�����_����1��h�Ώ����O୓H	�"�7�:�Ɓ��m�`�Ž[.��fE�U�lN��Hj���ڵ���Raqu��.��aup��0���rp�C��]d�¢�'�m]hm�(��I�ܞ8�+m�&�5#���P~���n#�#1;�|c�b�;��F:u ����9��(�Z�q_z�K�&�d�����k��Գwu�����2i�f}����Uu*���C�r3�48:�q��.�F��1�+�NG���4�t?�v��Z�M�2��or��8X.b��-��6�Jy�\!-�1r�I��bU�?9%kKc��Q�0�Ae�ܒ�凜"s�����#9�;91�ձ̍�:�Ĝ0鋀��1-J�{�rAO��*���Šz��IU�0�+��G�v���X*R3�^=���;t N����9"�b���>�E(��E�$b}%��+�m���%��W�LN)%��𷜘�c#�|"�^o�g�9����6��(�B��.���5��Z�/��z<!����6��Q�H�6^��j5ip2�L5�=��w���FK$�
D��W�IW_��T��<�ı�:ғ�B����4.���x���}eu�\��h)���vEjK�5�`�K��9]z�o�&+�RX��Ӻƺ8�p/J3�����i�%b�72�� �ɱ)<[Z�����ӧ��w,3�QG�$8���a��ׇ�B
����$*eB�OiL��R��w#��#�+�KV�%Z�5���r����N�����Ep���j����.ј0�Ӎl~>3�d�0�	`�U��3�g�L����$�0`E9٭������4�����9�{nηbwu���f��n6Ii�5��`,���?�0`�C��'����H�$k4�����N�]U}+ݺ9��s>�k�SÏ�`Q�b�s��{����`�-�DbR��E��zx�hȍ=��s�2�h���Ff7gFup��3�9��A ��*� ���%
����˚jcCK�=����ȯ�w?��'���#�㴘<0�e�>�η����� Sqt=dꐺ`^��Ϲ����N[���c�A�Ɩ��c-/sOFN�U��'�����DgV���ed�H�P�1}�BY�)=���'�r}�� �p
�a��Y�͜o\WqX�*�}5+y<�EL%]WEt;[��#&p�58s� +��pkǧ�M	 �^��+g�����2-fYПǅXY�sˀIFd����p���Ʒe�ן�a�qI�X����j��K0S8�.��ȇ��#���8} �r>'o�vK���ALp�vM<`Ȕ� �� � ��2�^{���Y��)wbR�{(N��P��&F�K>~��5-�/oI�0�K:�������C�L�<�dِ�;-�ؕTL6��p�� �- o�)Ќ%`�`�\Ԏ�cm^Z��`-N[�Xvt���)��՝�@���L�#0p} �~}"~5Ja9K5�΃0�#�~}Cޡ��y�K0� A��TN3F���)���ڥ9 &�k���t��� P��N P�]'�ԫ9ܙiWrb��k���a���%I�
:ʋ5].��^ؒ_}��8�8>��zRXM�M�e:ޡ�ך��3�9[z���M��Fe�`w��`������q�y�NR���*�T/�U<���Bl�r��'7UGc�U��ʦ����j�Hjl�:�Ѥ�g��v�L -�|� 7W����pq
�m�m�X�$ƾCNw������@X���#���ܡ�"G�a��R�4%�� �թJ��n�6�+�r?���Y��,w��KN-�r{\�M��L�t;�(mcu[u�j�k�a=�i�Ԏl�X��e�[C9��u�U ��QM�� Pr��C9?=ƓM�Dg�	�\̥�Rwԅ��* xc�k�Eʮw�8^|�����0�b�e?}(����-]�eR�p��jF>�>Љ0��e�s�/H�� �h�]đ����
Z䙛+Z#�i;�AM�<ٓX�&�.%��`G:'XYPXc��]�����!�ȝ��l���q9�"�Hn�ٴf�'��}vGu���5l�1�]j�0�I�=ʜy�^U��<=o �D��:}�mV��T��8S�
\�UF�%t��"��_<<�W`F�O��[�T�XrF����Y4zH���e��|V�N�e���L�Vp�I�hh��T}M�]�۔����H��2��;�fCb�1��h�4
F���xG����~��'% �N%��҆�{$b o�����G��.OP���?�����k�k/A��k�]�� ܹsGfx��T�&�� ��H�u]��ڊ_pGe�& �)�Y�G�v8�R�H��Ӧ1
�'�RZh�et�W�6pF� �E�|���X�	cdn@4�����ˏ$97+#u�w�%_�k�unqM�
剸}�W�TjI�����Vb$��WKu����,5N|:'y����}�y��B��|.���n�u�..r�駟�D}A�L��y���S�鵵5�ۚ�i�<qF�e����U��́B�qD����H�:VU2? 0�ۃ
.�*h����h��	��n��E�lA�� H���0�R���`}�L���#�򍧵?�L4P� +�*�� ���qw0�V��5��l��;d��nF���S)�8Z���p�@�awZ��g=/����-7��[��6@JES����pz���DAaw��������Ԁ��R�t9��.�`2�A+qT�}�nn�4J��٤҄�trb�W�8._�V�����	�k�r�`ST���,rU]�kw�F&Lwȫ����Y0^1��K��T.��s* �N$�/���ܾ�3��� �0�ƂdKMe�~o{��;�s 9�|+ك���1�$>���|����\�݁�o�HF{F�|��q�����d�C8�vJ�pn-��d����^� � i��T�a6+���� �fc<}=K�D�5����\U�e ٭-���D������r0��A>�*>k� g�K�� C#���K����4U�� Zr�3s��ՈS�!?��G��a1(�k`/�8�3`�Eٟ���8���$�ű��O{g�r�>Φ#(�Z����"��"�\GA�/�ao�u8�t*��{�nT� <�8U�&_�q����8S��9�H
̺�/J�Б�Ǌ38�=rJ$vk�}��եe�G�b���d�����
g���9��Qn�{��1μ��P�cdW�rp<'pL�t��a2Ti��,^)�y1,�q�	։}��ŅȞS�NU�%���Ʉ�39=�=8Y;c-#5�c PH�u$v�v����s��M$��L \m��tVz��Y��°�sXmwINc-1+�|M\ƺ���x�E'3�\RoVM���5cC����.��Pjv� Dt~s.W�h�"�'� �#�5��އ���Z�@<$-��S{��,amn�a��fe
�S�xZ�o�����iw9��/ƑI�k$+��D�ץ֙h�r��2�mVIv�`)���.�d<����@�H���2�@�iy�sl$����}�͜��Q���c�=v��>Y�x�=$� ����, ��+�<�"��Z:�rb�VGv�-[7n�V��J��<֚Yx��*��m�Pf��q�-�+ζ�kǾ�4P�<�4�˻Ѯ�HaͰ,/w� >�}U���%G{��d{�H������ ��*(|���*�5�[�iD�n`���`WZZb�F��������!��͈׹Rkh����)Q��hþj�~�;ߑ;�ޕ� ���zE.o��_���jM0�� 㩋�.��~ W̴ܾs�آ��c&��Tr����v�����}l��~�s�U+Q��!����fm����:>�S�|v�}�˳�0�=�y�/������߇�?�?q\��2����?����[�����޴ᱚ/��k0ƝH�'geyiU'��e��rb�$5)�c�<
��LQ��sQVV� r/��rvz*/�xEv�u�"�������|�+o�=zg�O��߆�����3����ܻ.Y8��I�X�˛[ fo������,u�r���e�b��=X���}0�����~��pd�Ͻ�3Bq��ܲ�Y곲�������蜮}0�i/�)��y�X��{��>��<}�z�Uܟnw�cN9���.��¢��r��o
Z-�.���4��X�ȁ�q�E[] ��mYZt�`�B��d}~��9��9��E�l���<#%nh \�5u �m:��� +%p0��6�V�k�����/h����L��&z[��ơ��8s�-�Z��XԞdS�Z��c��o " ق3d���� ��.à'cF����Nt0� �
���T��]�F6���h��R�&�Yl,7ӈY�;���;z�V��N�R< :����mB8௃�='w�����}uƌ�*0��xu�
L�#������Q2��-2Ȱ/�}0kt��q���N9qy8pQ�r�X]^z�*�9�@�u1#֎�b�hY���3�t~����|�����ǟ�q�U~e<i�(�1����F:����]�I'�pRVi���'���$��+>�X# X�F������2��#.��������v�u-�� �v��j�a���`�a�w<l�4�2�J�l�<n�X��%+�K*v[k4 ^�0�>Հ��,���ހK�ڍ�נ#]%����3�ݠ�;�g�8A*"�i�h20�Y�Zy������H�:v�°�)�������i �#9';x-C�4(��ܰY�z�=�35S�.����:�����Q�|V�pt���1g�;xO�S�V�Y6�i�d*�ڝ!{����U��Na�r8�Fm�1�L*�T��1m��7K9==�0���˱d�>E�m�ɂ���3\�$z��5k VV���b ����}�3�e�:|g>��/��>��yl!M)'&�3V-��Uǐuemt�r6IP~�Đ�AU���c��dCZk���޶6�(s ���� ���2�(�nd�!�tJZ��K��c�qjLMO��`��mY5�3�:�]b���y�p�Y��kh�z��n8py�
�w��'�@UM �a�+՜3���Qs��K�@�.�O����V-�gMX�0-1��0y�	ɍ2ڙN�:��d�4'U�^���p4��Nw�5�iJ��h3����N�+P�kͦ�W\���cs�6 \fA�Zc�9?���/��s��Er��~VN*�4�OR���ǜI��mI,��Av��6j�lӬP�4;�������bd9l� ��`n���%Q6$N����Z�ٮ�GfAƌ����/���8qF?��C�~������i#m'����}is�c�N[��YP��b��i�F����L�^��<a�]-�ٻ���Hl��ѩ���j������αV��cLY&�F����x�/�����<xx[#ơ�_f�W�~
rzx�peXa �W��Ǫ=�%V��TN&�YatG��u	��@�'�RQ}]ҩ�>?�}�i�Q���-�=<+��,[����P�|Q��ԅ���zx�o8���㻟�3��h�@��J�Ȕ��ayyUi)c9	�3�m	��5���yݏN{��*8��uȥ�M�8�֊'��a+2����? <���G���[壏?�/�+��T���aO���b�sx�l�'Ͽ�����v?���N��5�2 [ �b�NV���{(/K��Zr����>�;���wZ��$�sR*w�ބ�ǅ�;���L&�M������2�ݫ@��|�����,+���EF"5sx��r���`��oI�溏YB�¡�``"Kbqd��ל}��j�>�XY��#[�/���JN&=2�8ㄔ�)��er���*�b�Nk��N�F ��hl � dn� ���C�찘���ohz�F����A�\��)]o��� S�"Ι�8�]8���T���b� ��^wLk�Z�ဦ`Y�S����Z�E��Z��ӏ��3��'
���t�R�X��͢
�2�J{�n>�KSJ�a�2{�ݐ�y?�[�u,q�X`�JGu�$puF/��EZF��j��]���M,�Tj�z}~�������փ j�õ[Y���4���5
���lT`4��X������
��ryuN���K�[ d�K]���Qc��g0`���\��E�XV��b�~=m����C�8h7]p|x�Ar��X�:��i��ˑ�	 +�*�S؁8z:��a���?;�O>xGfXPvK�����R��B�&n���Ơ��o�p㢳�ެ�����4ᐛ��d�:P�u��V�vnX.�J�ߨ��lVj�@"XGi����SV�Q��#q�]�I�<��C�;�F�Y���h�J���s2b��]r,�i�I5֫]�4�>��]��Ms��\�3�K:G٧��3'Z�cs�h�k�ɱ��Y]t�|�t��ރ]i5pDpN�H�M�kr�'	��%��W���M���6���a�?���ȍ*�?R�]����A�ʮ� ����pJ��`��]H�3�{S��:��Y�lq�Դ5������G�A'�wSG�~a����&��ޮF�= ���d�.�}��p��L/��C�X��v�u$���Np�av�e�=cP#^I��H�%�� ��*��-1�&�_TAH��p"�Y[�X�?�������5l�ƼR�}4h��i5KDd�˂�����t[mM��?�����9�=!�)����0��FT��B�X�
�t���QW�ɸ+�K�-t��`Z�i��Z�S�3�@v���V1��p�W��A3��Y�r�[2n�J{E}H�}j����먲z{ 2�U�F6���MM�2Kd�pR�IS��c<:�(��Ĩ֕���M����>#�%;���&'��-C��f�1օ`p�3�n#�@��D�&�Z�����0:��}k4�[���1��{w��y뭯j�B���d��j��Y--������78!��^Á�Mqf4���g�T���j�m������J��� M����)������?���%���dmuQ.`ְ_����uL' E�f��27#-j��:0�i_�./�'�+i="k�N�K�~�z�2l�EU)J���E���G�n�-��~�� L	#rv��ϔ��� ٨�����tJU#��şJiz�����vͥeY�mc#k/9��gffV#��>ش����<�\3����EN��6p�^~�۰���W��ZJP�洣<}^�߫*в $�b�fF	������Rζ �R�|y]�Ų,-q�$ִޖ	�i���_�/���Ŏu��).% �Dr"W7.K����jf������Ae�:�A�^�) aM�ݶ*i_�#k
�y/� hO�<�3L������2FU�ntz�S��uʐ�cVp=������G
W�'���&�h�t�rr6�DS{p�!�]�Q84��ϥ�(����0��2Xذ����,a�C�a�7�4�����`�)!:`:]Ԫ7�A�dLd>6#vl4# `7v�MLZ��w��m��ܼx��%��;%��U�YBvf�l�zXd�x��:L(v�:( �dܠ�'�z�~�i\�8��<>OK*�S��X�S�c�=`��8��,l��lR�'���q�g*J�����p�0^Le�sKl�U��[=�.�ԛ���X"�
F�� �l2!h�� �"�C�U�i��Vn����]��K�n�ƍ�NB,�/U�ؗ�$C�f[��޹���|�)YҴ��{V� ��}qbO}lQaV��=V�w��iǥ��������)�c�N�(�\�*KP��,��Ԯ=��%��|Fu8@J��b�G�>��?6�֋1��тf��:G��� � �K�Ȣ~p0F���8�F��_
�2�wX��) 8��,ZmM����:LO׌t�.-Jb��E���D�Eu���Y�PZ��2=�7��j�< ��2�9���մ���'Ӗ`0*6�kt2��3k� �'�O�.�N�EMC�K������'|:���d:f*�� oG�����
���Ϝ\���Üc��]iu]X�9����L?�XQ��5z��)x����QD���Z+iM��hbůA>L�e7�Qϣ����+i���,��96X첲�({X�>� N'�P��I��4YhGZw����H`-����Bg]3�f2Z�!ic ���jAoPm���~ڸRam��#.k@S����	@v���!����p�������i#�f ՚>Fm��� ]��Q�$�&H>c9��������vG����M�q��ćJ|��q����Q[Z�.�����hQ�`��Ԓ4lA����'3� ײ���$�t��D�ƴ,Ϻł5\[��Dا���ή���`����0=�O�A��T�=/��$a����3��"����`W�5��QK�V_Ё��i�H*{�rT���$+[� ���6�1h6�~����֍��8S5�־�Ө#M.  �v�]�}1���aZ���-t�ݧu�N��;��Fe29Yݸ�u־pR2�����&��i���:����c��e8�A{O�55�sF ��xd&Ӯ�J��3٭$��������u�
HjR��$9Y<�	�t�9�;BP�q;�Z����TJg �69�"�ٙ�d�Y��:l�Kӭ�����cw�T�A���=��9@XY��A�27����Ǐ%	�4��ϻ{t4�R��b��r5'��:��h�DG�]�����J&����]7HC6:�sT��u��+�͎�!v��1��J1�_�M�\1�ʉ&��_�D����?��%�3k<��_���|��etʘ��ю���Fڦ��G2??��o��#� ��iriS�f�U�pK�ڃ]�k2��s��buƥ=l��ڈ���?��bH�\��.p���j��&��		���i)��f0�b5�$�!��1���'�l�m�i��-��!،z��kn����j>oP�L�tb��T
:���ا��O��B�a�6"�i�|��\F�����ד� �`ٙ�m�YiV�rycF��(8qk�΂N��@�^��c �[�a�Cވ�cvj��נ09tm�d1:+�pLǻu,�Ͻ�m&�i��P�?.ֹ|��k�3����-�3K`q�i*���ό��\^�V1u�g$�bM��U���;+6���cF5[��H�� ��Ӑ=;���Mf�!�f�,�H��W�_��~zW.m�J�5�����-�u��s��Y���+��9	L��-��[Y�SYcE��|peH���4й�mvtN�+y��h'��aV=�|�L� :10�. � md�S[����y�TNq����e\# SCe��F�鬩�5[�P��W$��4��$�j!#�SS�~��j���f��eŎO:*,��
�:��=���Z[�8ńavU�o,W0�2��(���N̨�:�\A#�t	��˦���t1B������w�	�H�[b�-������;��1�(a&p����`XW�N���D���%�(�u�V8��;$�������+�!xP7:T�� ���t�dٽ�jSM`L0���5�qǅaox��:�g@P�0��ڽ�I�?|O��y�e3OE�eY'���Y�r����+��Q�s,d���b�6����jc1�:�:��,����~o�{G�E�Q�U�`vhʒ2SC�&m1[�z/N��:���3�Y8���` L0���V�9�d4�5���5�a{�Xo7��=�4��`Л���.р�)p ���5m��1ݷ@ҚbΊ��޺3��_0`\��{)���Y��E�~�g��ʊ����ɣ�>� Ì���;�Y;K�4J�������y9��\|z�HÕ����b]����I-�:���Ʃ�WM \8���
�Ɯ��Ӓ�a�$ˋKb���Q��#� ��ގ�2�l^y����`�]�&��L��=��%�����+�[ e}���AR�})��ԕi�N�����N��^Tj��ܓ!�N���J���� �����nU�gO�EB�t{�������Z�*f �No"E��XЪ(�</\/�Rt� � �4�.��^���Ď�46���Lm��ݼv�ϯn��ǂFgW��s������S�7#<�]��+N����F�y����05LE�)v��q<����y�y�Fz(�V�7u�����[>?#��<s]�fx��	��ZFu~q&��d9����zE�'��)���k-g42���\Q���SR�A��i $ð�߿��LXkL�p(&+++�Z�iZ*�]Q�Ø4��qB@�����X��
n߽'�s�2��i���$a��99>=Q����'���LF�VW��ۚ�O�N�f7���kf �݌\��'��;0c���{WV�gp�g��O~-�� �<��HN�g:)���`k--�}�@r�`�����N$3y`�q9=:xv�q����[��\��T��(�X@}'�%Wօ�pM����UƤ�����a1�q|��y��Ak����Sm��٠V]�r��J��}�K�6���Ǐw�&�&� ���ѳ�y�6ц��m���b��b$��l8d:��7
G�y±&F-��'�ZG����9G��0��c�y��-��rZ��6#yعXL��E�C���������H�:7��T�q�� ���\�p��^� �fF�nw���gS  �*�;�w5��6em6!>z_f�~yy��GT
m�9��c1�y<VUH�k6�0r���
��h�4�J&�SԚ4'~��MX�A#�#�c|��j��(6ǰ���8/�uǇ�z�Y�����v�9����jZ%U��`rv�1U��Y2
'�y� ��qD� ��9�Q�d���x)�~�5���C�d0��?����Q�������L���5x��HDm�w����;?:�d|@��5m8�f�i*|�*�4���`K�:�{i9.��9�� ��_}c�`����alǤd�u��Uk�X�����`��QW�
	��0��:`�N����iѮC�Wl`��#�)W�+���p�� R�ƣ2�:�	�ɴ�R���E���aY/Wg�J< ��#�w��]�s����\S�����p�;����v`�F�	s��²[�A3���9���
�]e�n'����=Q �/���3Ri6U���\3�V{l��-*���N�N��8���^�jj�	�J]�A=-;Onc�@��D��?=<��Q}2J��iw��+���pguM���D\ k�i��$���ڂS� �:_�k�ւp#�����f�Y8���G�9cT����I��=�\�f�'�l=��Z��b�������x"�
`8䴐~����)<�ɩ���ܨ��ub�!#mF�u�x>����Y�s�h6�,;��@T>v� ��Fb��K�Z�{3*U�H�_� 2��!p'=��x���9�i�����.Jw�����$�`�D`Y�.�H�~*�@�1�c��j�B�g#���<�#v@ɕ	�%�� ZfBp�� ���>�W����%�����'8�}������vR��2�C őov��J���n�+� SeF����kb4{� v999x"/�p�z�-gY����꼔`OkEj���z�^bo�D�]�x� [&7l`��2�S�es��W���&D�Sg��-�pOݰ˅�j�Y�c M�ׁQ��u�$ \tE�u\�AǸ5�` 2�p��f02(����x��,�lJ���HB��_$�����i�C緐�k4��j��Ǐ4J��s�fR���7_������69Rf�v�t�?������:H�G��������{���F�^x�y��?�#�DC
ON��5�l!i��v���BA�ֺ�)�L��$�6�4�U�����;�߸/�A0�L	�������=D<x���5��N�`fgU��rK*�H5����Y��]af�@��֦�{櫯�!���f�*�M�X��@��Z���	��B!��{�5�̧g��a�N4��#ׂ � �M�|�@ �ޒ�E�ӏ5xs��e��3�[^Y��(�N4JG��;�2�HT{��@6�/I�c��3J�4ֆ#3/�{>�;�-Ij��%vhðԧ�o�D�a��9���B�"�B�00Ǿu�=�.��jR�s"˫�diiI>��6��A}/K��|�P�!�u��`8!g�ǪHB�^�^�v��j�MA���~Z&3Rm3��B�8���=0�ݨF��7qԎr�س�'0��Z`g6��<.���pH��L�sL����m0_�p��>�3	�a�����Z��l4" #1�o�+�#�rN*��K��vGY�2b,C���ܚK�m�#W���vU��5o���0��Lf�s��c����4���#�XTdb�VϨ#��dX|W�c͍��b�p��^�Tj� v�0p���v�����[%��	RSG����=8��@kx��rp��`4Ģ�l>@+|�_�>��RL���.���؜_/D�h���Ѻ�"`����e¡+K�"z؆ u��>+# l'`�k���X�����l�xZ)�9=(V av��l.�@��l#c@�֤��G�sR�ݳ�4�&�9r�嗥;0I����Pe%���~(c@0Έ�`������hԻb�`Z�F�Ρ� �a���Zwȼ�y�:D8<�]��fR�l�p.� �mib��Z��u��Z��l�ӡк����m����([&, >d���4�v���[6Bqڎ�b
��(l�2c5���d��{��t^��T��X�i����jԕ�X;���]:}�>�d?W�z�>���`� �2CԻ�x�o��9���|ϛ���F��!�W�.#�QU:��6�P�1��	rp&�^X�?����-���.naz8;Mq�<������ ���z��h�4q;�tN�զ�Eg�'
�t�p�N�o)אj��nv	��aC�Uq�n���s��Qr��/�t��"�ͳo`�v`�Hh�ӒT���Qӻ~��u)�Q(��,ʝ;���F�
';�����ƴi�q��Pt߁����x�� �fQ��q�p�f�8�Xʢ깕�Y��÷%��r�ѹ�a����e58���l='�3�- A�k���.K����J��L������^�$.�TC�=�˥���ǘ����<SG��h�t���	�����T3=���. B�ek�ړ"]v�����58�FC�â�H�n��Nj��7Pr�g�btI43i�;dјXq�C��j�q�m4�5� 	��[mvaw�sp��a7�=;�ic�{df��C��k���N��jp�s\-x7�c�.��*�v6��̢���ce�tN�e���fd�#���Q�vp�K�8���Ig��lK<9#�\U��R�dU�-Y�E����UM�NL�n~W^y�%y�g5r�uy@�Dv�XJ�=�t��c%��l���Hߝ��e��Aj?�^�w�G��λokĶ�n�����0�L�Z��}�h�6ߏQ';�e�ԇm���0��	���tD`A'`1"h�}d�6���?L�����i�_��c7�ΦP�*Co�/:�b49��+�bıV� �U��|=�U
a��Y��c�������`@�4�ͦ.��c��ڵkZ��x&8�6���9� ��jUf������k��I��2֊
Gk��t��LR�s�2�q����@B�7��U�֗��[��L�f;������<���,��e;�>7u;�*ֿ+ONp���z��%��N�N����,$�+�w�ܓ��T���g����S1���pQ�&����JXM�CxWJ�Q��{�u��&�]g�M��ٙ���$(��v2����ᶄ u̘?~�I��ߪz��s������1��,S�G������&-�e�N���T	p��YC&۠�ư3��\V�T����@�P.��CjV�JE��x�p��b�$ҬU���C U �|�9�2\I�_ �i���^��xh��9�qŁ��tk���uɌ�2��򅤋��IdD��,�!�9�X�	��u�$��KQ겴������yT�Bbk��d��9��=PSʪ �#lÀ��nM����-���TkHhaQ��x�I��k� smi��&ޟ)��X�#>�PrV��̷�}�>>g�p,�FV� �UF0��X.on�ɸ�UNK%} &��!�V�
���Ƃ�������0��E�	��jp���?�Ѯs�N�R�����h�0
uZ����{��J����>p�Y�8$8jJ�p����`DjX'E|m8�����g���#\�y� �JR����ڥ儖A��^��P���]'�,-�H>s&���;�����T���T�y5�B�)˄�M�J�m���|XZnֲ�0�G��a:�4-��x8�c��9R	x�(�xHG/u�mv�խ�����w�PȮQ�G�#��EE��*U�_ ��/SM�Z�U�?��_��QQ�w���
m@oV6/�$/�����������H�ÿ���[���|��l����l^�.���d-pxn�7�]�.�4u�{0��y��CQWvq��]�n��A�Q���~T��GB��JXs�uv9A�n<Ǻ<V���2�|Q��ߑ��M8�+p2u	gq& F{8����nu\K�k X���'�w95�]���歯���ޓ_~�_�VĤ5Itn?/�����!�P�Q�[o�}�ͬ�;����>~�H�,�`$�|�S����!��D^������U�Јኘ	i��r��6pK�`c��q�}�]|@[=#n �����[��8���U@��Tƃ$)_9�H`��3�Q���ee��u��+�z8�9�53�Ҩ$&[����0� ���
�&�K�Y�;-h��R-�Μ/��\�s��� ��R��%�f��W�}��*1ʔ>��7�Ԏ�>'�_�!�1��3����I�`��_� �&�9)�Y� ���q���Q�5�S�� 8 (-��A�9.�N����Й�,[�|��u������<���qV;-���������<@�#�׬��� ^1�h�������~}��W���eM$��3M�R֫ T�ͼr���a���w��k�)HdƇc#]<>>�·n�`��{�r Θ�ʊ��0��8�]�f��.�!싁J��i��́sȮ�!lk!Y���>���n:���YL G?�p��YF���=U���]��ӲRٌVC̬�7�E�B��	�S�=�h��X����_ʤ0=�����X�kd��(�����BI{1��!���Fh} D��4��W�n6<g*������;wv9� �  ����R9O��ɡ�o��
���+OkgO���To�G� ҦZ�ɔ���`](�'jU��4�ן?>ģj�|&�D"^}ߘ)��M$�����A)!�$p�ז���| ^_T������e���%��q&�(,~"+k�:��D��	V�G\��ZP���i--��ᲒX�p����(4�f��@��v��쀋̓���qߤuN,�g=��dlQ�<���IS�������3�#$e�	�ـA]3��z��52�fK��K/ܐ�xT���VjVdd5hmR{�L��aj���n��3`G�O5˵��NӚ�3r�Z�h��{ǋ��!e����V�[C�`@kN. *����<G �5�?c�b�D��I2-��w�r���K����x_ʬO��Y,=��?��0/�9�Ɯ�� Kv��Rl�4m6�s��H;��3Q5�|g �3���ʦ<����rUך_�XTX���G��5eg��O8� f�
E���9/J�Vǀ=�ao(�I�JL@)%}p��!'`CA�<�@�5]�E����7a>5�W��7�u4�NQϼaZ�p�{��5�6����VY\����V��� o��17Aנ-�|JF AF8! ����Z���^�E�����Ns5I�^��ô��O l�8������p/#_~�U�*.�H*80�9J@h��;�ޓ\�1 2E�Y���9��Y�N�'�l���P��a}6�p�١ڤt�	�6�Q�nS�$6�R� ���И;5[���P��y�&JYa�n�� ,�~����!��;��:VNʊ��pG�6Չ���g�o&� &�S� ���ob�p�Ay��ߖ�O�;ܟ����������<���ߐ�����0o��3���|K���r|����ϝ�ޒp�Y��N�n��ҝ�]�W/���%�?ޓ>x_k�輒s��w�<OI��O�C�	����i���+���ZJ���8_ ���Gf���w�w�W��{�w�����׾�η�!�;�N<y��B>�~ !G��\��"�ˣ��\RB�n���ev��hCS�Ȫ�]aY��e � eK'�L�6��P����7S��Z P*�2je%���u��W$�q&�E�$���-���xg�H x;s���nbӋ6��ri�Y����pL]-�'1���w��pq%.�~Y:]6����yS�����W@"O`��ƞ��wna]�5��_�i	���_,Դ6��5�����K�
��X��Q-[�����;�w�_�0o�w���� ���җd�d�3ѦN���ܒ�� \#b�ΐ��.	:�M�՛J��� �����-=ш #��ҙ6���T! <����@Ч�h�}�@M���%�1�n�D�&�R����%E7�{C�/z�N��1��?�gn\����l�,oi��Z)hѾ�h�f+6111D{����oJl+���ssKj���2��5`���/���>ld� �k�(cd�5űXH텎J����*�܂�����������m	�v�E�	�c�}�6��-���Q=>����r�Z�¨g�c��ftpeu^��� ��������a
���d}]��P�����V��0@Ù��?V����;ֈ0�L�=FYg����{ݖ�>�//�xU�#n����D�k�|��/�gF2�0?U^PMǪ~6�}�sanA>|$=�8�� ?}����3Z�+�Շ�}r����Ѵ�Ť����(�˱�+�*F�;��-繜d _�r4O�_	6r�/���'<��G���y�_���;+[��ni�˥���doqnNSɬ	=>8�X$.N���=�2��lL�)���N���UJ�SN�Έ�O@:����n�u�a9�z|A�O�N$�ܳA,��FA���l�Fu�cw�#u
F��6��Z"��*-0��T�)LOGr��K�3��[自U�����̂d/���� Q7d)9'E�6{�Z%��2�ccF�>�4Y#^�v�Y�,Wsb	YZ�V���p�I/��" ;Aq�ul�8��2��7�@[m�l_�U:�c��Sl8�N�M����u�Fn �/� Fp"� �4�<�r��P��j���y��YAe[M^_Q-�j� �s&�0$�u��`�8,ԍ2�%���o<�Jܷ$g�b[�i��lk��"�p`a��2j��,0",�g1.���s�!eLb&,�t
k���)�tIA�㇟�s�p���SD�ric,0���=�^{���N��$tv�3H&���6�M ���Tف!�E���!�n\�''���j��A8�N���#�(��zEV�}�Ka|^_��/�Ċ��`�)KAB�9kȽ����I.�I�eМ9�'K���3��G�gJ�R�h (W�YR-���Y�z;�3X���������Q&%E�/�=ꀍ�jZ[4�!�6�a��b]5�(�df�+#�BmK��fd����M9>v;�1a�#�6��;
 �n���0�y�u81�+��#�#& �~ ���&�hB����J,�[/�(V
�Z`L�6�[}N�&�>�-�qWn���dse9||��	 B�������6�} �ȟ�>,���LA\�k1�y��_�����n�&��_� W���qS6�� �ߔ��9��c�� ��1��_��[W��pl^.��mF��CZM�������%�ZZ ����~�
�RF�k�x�̭�I�t._��ߓ뗾,�tNS�'Q���˛_��l\}�I��s�?���c=*�[ω�1�����%}�v���7_�@,!��9��z |!�]g�.�A� S��MJ��	�W��XXZ=���)>���]�Nŝ����l��%=j�g&!%�����T�PZ�Ėn�B�!_���΃m�����ɖ��z5(^k@� v��b� �܇���֭2�Tm�����9�qeC&8G�l
NۦSH����-�bNf���Z�7�%1L��#3��<�D�8R�m�ȭsz'���ZlC��Lif�9����EIu����v �(U�W�����Q�Jt�c�v��`y�FC�j�=8�4���(`v��q��$�aF(� ( �v_HL�ɉA iV�wz*��a��p**�����*,��"pt��bͤ�C{�RFꮲm8`�^�����KSy,����<8%��׾.��H
 �.�'�
���u�'r���-Z[��	;�{m�u�%MI��^��-�P��5�/ߺ)��ym��{�rqz؇�Z�HW��3S�k�T��Qu���jf��
Lh*���_�ղf>Fc��mZ[K{C�T�Ţ�N�r�Th):��\���KWk���9-�r����-؃ֺ���s����n�
$�(�@��[�����LS�,02F�P P�8�ͭ-}��Uĝ��Hj��9��w�G��㰇�:��\n>sU͜�GF�Pb���K�6��`𗹸�;̙[��w���d�	��:�5�&;�	�U�A�ڪ����U}Ȅ��'��g�:��
�mAR���=�H:䅛�������g
�2����b�NV*����/_��ϗ3z^Y�y@<�rpr(+�Tdí�8�|�aZ���0�cN�aM7}z{��g����o�,E�p�@�)�^ߠ��w��.ԉ��M�y��m��L��@�f�i�V�w�2#F朸�df�lN����b�8>;յK�e���D��*�0em3�48�R\�xQ	 ����G�"�ق\����5	z�`l!��)Q��jmWK;ج:���;�ab����<.C�[�X*�ylR�� ��DF�,�鄗��8P�RW̺K�y��L=���(�T�,� D�ؒ��O4�c�sF�8�0zK���"ed����M�������Od���,���Q��h�����`� m>�{��ܳ���TV����G$�e4�L��#B�
�����y�p��s_G�l���T������+w����l��vڒ����^���Ei�/H�Rսay��jT�Fd~>en
������	4ZMc���ʶ .F�`e 3��ߗnl���)a��Q�"�^@�?ݖP$ {'G�{��/�w��{r�)p���[ߐ{(�^�9Hi]� ��Ύ|�g�ai'#k�\�����k�Wϖa� �W��p���eu��Y�惑��d�u�f EE�kY�ʨ��k��Pn�`Չ,��<��]%\�͚�X��j��ӂ�-*m���<��W�łD�~K��1G�ʸGc��98�!ȃY~��}����*V��cy�_����۱��?�23�%��=0����A�������P����#q6� d~��6�q N�+�z�]y��Uzi�g��T�?�H:�00H�W���geg�1 N@��o�B�bQkco�v��?���H���QL�)��x�_����
 ��߅<{㖜������������ x+�P����d�99��G;��n9>���~w{ �X˾|��#Y��i�3��X�<�;;�r|��� ��pʊ[~��GZ@��PQ�a�S8�f�-�Ӛ�?=�9�W�������ى��%��#%e��M�uS��g�R�H�ۗw���$�n�,��W<��6�&����j��� u!v+�:��Ǐ���kCN���Y�ǩ��ϯK�6H�ꅜ����Hv�p�'~��ݪ�h��|�����nUm�FM4���rvr��B��h��#�Qi��p�&O�ߖ��}g�%'ǔVqJĆ�1�G��H�K��$��E�~������ը��9��4�=h��m��$ [psRG���*4?��@J�R)]�t;P[���<n�}#h��l��V��k_�����`_;�%���L����N��ߚ�Plz�Þ�>Zpw�O��ח����N��>A�H�U�>���/��K%��12t��D���rM;�)��n���UJ��@��a� ]��< �l�@`�H�QԲ�2�x�p&>�)Fv=���G�>��fØ����u:��nf�<!|�!l��7P�H����ҕ�*	� Q�I&����tKr&.=�����T*�2n��{�Wp�������_������%���׿ĳM���ohT���lV����4�^�}y�����>�+�.��k�P>��C�A�tJ�`���֭[���s7_�F�)`�;O�2���}9<K�lئٹH���ݩ�O(�#c���`�U+�z�}Jߔ����4�y�ϰ){�5:j��b}K r�')	��l^�_̩3��qo&Z�fu�$�L�?��q��U�6�MC�:x�*YU�=غvI<Ҕ��Y�{�̠�u�x�z�d|K���f� ��� �I�8�?9�j�.��,�~G�1�S.U+=������B��Xsbb��0V=)�É���c:$,�p�@�C�T���t\��ڗn ��T��lP�cO �qa;͊x �J܏�H�`����U��胓�1�ʭ#�4��i`{0���.K��F������9m����T�����p9��х��+���&x�n!�A&��k6t���&`��@�n,O� ��ځ��N�S;]����U'��4U�ǥ�gt�B���رH���7$@{��\>��7��o�#������,��gߔ3�Y�6��"��v]V
<��e�����K;��%�{'��葄�!8�lݸ�� R,�����SE������f&��#��=���]�!�@6[ �������� `��p\Qq%=�>���3"qօD��$��1@^��}�|�
΁���bT�Eo8m����Ol��؋��N7:��!!��>�z�%���[
�3xEם
`B3pp�%�ʫW��?������䏾��-ܒ������/���v:�h�	cށaؒ�`eFN!��%��ku�d�N��J��=LC�lX-t��X��͊3LY�+�g�ic�ꨙ4]4rME�����gz�)�0�yg�V ��A������12�aE�h��,���2��}G�qj��R�G ����Z�DF`�Q?��i����T��˰����@�&�}�F����k�P0����	��d.r���k�<���0R�qy��C��ܾ�]��2
�S����_j���%�(�ѾԷqG��;�g�ʤUȗ$��,�����ӑ���8]���H8!���K�W#{��b0�����?�H�{{G߇F��siCW�P����sի�xo��0���C���]�!8�\m:��3��C�sb*&	��c����ӓ�
3 /�Zwd�{ �`�G8�^)�b�d1F�,��`k����[u}���/m�l���?�9�*��Zh����̂l1�A�D�N� �2�$�wk����oI������+r�+����bĞ��ץWJ� {�5z�����(�?�P���=鏕�x"K Pɞ>��,NO@���~8R{o�����fϢ�Y�]�0eKkA�[�M�Z8b�ɮ��a�r��^&n��9q
�G:���<�;cƹ�Il� 9�>������L���.�䢘mq:��6�/��/���	�:��msJ��r#3	��1��"6�h���G�F�-���R~��G��D!���;�_)�������Ձ���,�gL�oߖ�'ߕk��j=�[��EA�n�g�X`�Ւ}�cF�`�:�Ɲ<�Y��y����/�(oEq������M���Աo�x �*(?��ϱ�ci5˸�~�,$��6����懲˗ ���P��pv��9��bш|N�B0����-��v&���[���Qkv�U�6�YM��� ���!����)3 �̒x}98ܓ�ԥi����<����K������<z�0n�/4�N������ͩ0� �ly�wt�
���⊄gr��]���0�ɩS����>��w���s%U.�ӥ�8��_
��ZJ�́��Jr>�s���(HriN��]X�R­B�l`u���pD���p�	:Ov�e~a]
�
ΎYf�٣m�t�,�g>���w�.��]�_�Tq�;���$N�ۣ��k��4��N��v�������֦�\�HFFO�qK"֌�����H�r^��8�̙�t�3��oNX�+�oo$i���=yߙ��YY�]���1��s�f/�,��J�/^!$�l0���0&�!� ˄0ˁ���J�;�evgvfw���鞾������ά��N?��U��^"�&:���/���{�����
�,�$�/�F��oB=~�E�TG��r�X6�Q��E�Mϭ���\��)4,���g�\(Y����Z�4�/ki���r(����Q�J�P�Ӂ�ٛ.W��X�WGpx��q�����*��8���@S�3j�Xy�1ܼy�8��kOP���c��<.����|֔��<��_]��K�p�ipBQ��t_�*���u:F�l�=Z�\v�:�t���oݏ�^������짿���|	k�w�Q`vq���z�����q����/<�g��"�y���l͓���?�
WVx�n�M��+_�
=�uK1�8��g^���N	п�ҧ��N�R�2�*�6�({�K�~{�1#���$L��v��@���?�m@B���n����U�!�9u���j���M4=*�V��"����]4�L�A�L[]^���~��5�̀;q	���&��x��6��g����
����oc��g��_�=�4�s�$�4��^���;W?F�Y݉{YK��y���|N*��?a����IR�Uu+"j�Jæ@H޽F����dF������UP4���y�F�,G�(������?��Z�tZ�|��֚�8,�+�	����F0~%F�ܡ�y87�5��8xz���"[޲Hg���k��Ɍ0��?x���*@���)��j�4��s��_�
f����Y��g�������:|�I��<�����6brz���Č&���[V�;���K��mnd�?Rw#���9x��K�->YB�gA�Z�0��"���8��(X�Rb�����q3T���g�yڨ�*Mu8��a�5��ź��V;W�:?��Q_�g���<��r��-���*����hQ�U�;M�3��`O��2!/r�HLL��;7���܁F&��K_���˕��7��E���S�V	��#:��9�#�0�E�V��zsf�����/Q��������D?^���p��o�^������H��OL�<��q�x�`��%�H��)�G�C@�ʵb�k��:\��J���#��g�<��@\s�	���Cf���GH σ�~�4�j����-|NM�7��(�<���i����>�x����O��Ôˠ�ms���i���=���M�#A���H�K�d:�\l*+E�����B��A�����_P����!�T�LK�ѨR|+���5]�}*���Y��=��n�y��]��&��J�Iޔ����"����4㓥U�:LƴQ��89{��猘������̝����櫚	���.`���	�Ɔ��H�9:U"��p}#���$'��,��Mk�T'rC)dM��h@�)Q��v~Tw��ܪM�*�	U�|��YS����9�ݩ.�a9��4���ի֭]��H�S���M��0C`����ޱh<�m���ݻ�0!�urr�P\������j�\2?�hQG��ݿ?����K���})�kG��,AϤE���M�}�>�k�J.���������� M:=�t�.؈٢5d��@D�HP5�*1����c�^����R���@ؚ���%��l�h�W\���-qob��I�W����9tjK��*_�1�[ow�O8ئ��Y�Ï	2��[Ҝ �6��.{~98��J۫\���Ӡ�����2��]�UUC����)'�����ݾ�X9�O3�O��w:�N4v���|�MoQ�s#�VN��3c�y�!i��j��*�b�W�^�A.�a�tj�	�"hQjVM*��"p����ϛׯ��y
nAT�j�*(T��T4w�a�f��Gz��z_��&fy��C����k����t�.-}H�VG[��H5~�L�bAO�BO1��\³��2�(��`�J�mC�J��C�zL�B��)%�'	Z�w��?9v�|��+O�P���{�U��=�����?�V>�AzL�9��$�!`�\��Sg���n]�FE���h4�2V�-�J�t_�����_�&F�q��%���P�O�^��؅�7�T��!��˦Hd�U�0;g�w�A9�[K|͢5*��?� }��V����������K��䩆R��4��Up,�rq;u�d�5�C��r�p������n��^�J'-z���P��a��1s0z������c�{t��}�ݹG����*�X��p�F��qh��������X�o�������1��#�eO����ZQ�F.�赟�^\:΢:UW�Fl���'���{-�M�q����"�2N��Շ��&Z�\�@�`Ǧ����
:eF;�s�K��(%�Z�@���.6hxW�v��8Of�� ��H��(��`ǰJct7��Ք�����}: C�ߩ��404l]��Q@(U1<:f����}UsZE��3�������Q8n*2
�Z�,�_�X�<��eE�h/���MM��9�i�Kϧ^14yUl/�=�#b��ON����Ѵ:��5��$8_X����9aɴ�/���JA�0j2����M5M�X���]�#p�h��.�y��gH�<3����Q7���*�Y�ް�R�����F������t���	����N�x�1��Cg�J����
��H*c��>���~���m��t��0�]=x�������2�����]\�<F�����x�S� I�t�c��]$��e1��k�[X��3ǆ)��46���>��ģ��t�g�;�^l��YJ-�H!a=�_��cp)��ԋ1#��O#C������A���K9ר�ϟ���v!��c�u��,�*|�Q*���œ���V�[���ߓA&�8@]g��u�J�2H���@AQ�~l�~>��]�
D�	<~1Bxm̧�r�襚q��>u�.���3�,U��>(�XiB��X$��v��QQ���4����/�Ep�������ƭE��[��7,%,����`��z�@��O`pe�i܅F�\J��R�}<+��|����r��j��ܣs�J�}��S4�Iܒ�<G� u�a���I5:�6S��6'���	�V�>| �ۜ=�m1�l��XS�tͽ{�8�)E�jM�GCv���28n�>~bΉ&��7v�#\���9�:G���c6�����c�������+��8�A�z>c�q��^y��'���*|󏾇t�Ǧ0�jM�^]�\J�<u�ؕ�l��F�E��3���(I�����.?�"n��/=� �m�z� �hv�I�S}V�"ڣr���̈9�j-p���f��t�2)� _�c-�����J�Q��山�iI=�����i�{[�@Z3ē��Y�����h�|�צ^�cD���b����g���&j��N����qk�\�(75�x���Y6D���:���M#}Õf�S���B��Z�:�j�墀k�G�B�Q�\(dC��P����\����Jͦ�!	��V�>��� W=G�E2�)n����U�5��w1H N����nOl�T�*ju�]F��	���-�����!�Rq��|��E��[t愢^\l���E��EMr  �����@��o��,g�+��A�j��4�
���)�5u�&�� ��"k�rXX]���E�&��VsX'�X7����jk{-��y�Cq���,�_{c�~�%M��٘+q��2���)�����c\�*٢Em��`b�qC�#��6W9����:mԸ&J�G��5�/KPP�V�����ݳ�-c+��+��8,*v:�|69E�K�8s�V�H��Pfqm�g)݃��f�j��@�u���� �G�vkc��q_�@C�H �5C��}���O�ݫ�Rc��էEH���]�o���v�׳�sg/r�THn|���Uষ;����������.Y�F��juyψ�c�寎''���n���5��6У��8e�LUh9
�6����@�y�����LM�P�w�k�ȸ��j|_��t�$�:xH���nd	N��)B����Q�7�.Ao/V��{�(�D�S�u��}��/�P����=�|T^W� �<z�_�����=������<H.���ӗ��5�W{/�(7;��������G�wxx�8�d����{E���ϔ6�qa�#]K����D����:�����?��9j>�k��HNuM];G�H);]G2(�\�,y3#(>��gճ�y�Z�� �f�+�<21�*׷!b�|�[�`bc�a]���R]�mn�ཱུ�`t���H�XG��||t/?K_.��S��BG����\y�y�ݿ�w��7����3�����/�E+���_�?�����p�8�����7ަ��㵕E�B�E���A�D�os��lr��p@���g�hqm��s����,�|j5@<�s����d{�� �����
W�{st�n�F}$ �N�6�1�})��ء����"A�dph̢{j�r�vS�ܺvݺY��}����m���yո4�M,.=@�`0�mM@Sό��#�?��������Z�C5�"*G�\�<���8}�ܾ���+��+!����z#�[o��A���Ċ��	*|>����ns
FGΙ�3�}��l��u���C�M�|��(��̅�h�[�-Z���&�T�K8�;˿9���զ��ղ�n��ش�H�]tV��m������T]u�X��&�h"��Nx�Ɓ��EiSP�
�W��NG���@���1"zW+`�ܥl�"�r�S�N�:F5�jB�k�´��z���;M��Ϯf�sg�`{gݦo�U+%[�
�����}lgptd��t4���;MkT]���-����<l/Ϯ�%�G@��|��N�I�yV'���ʭ-���+W��UM��ŉ���o�6]$K�ٿ����'�-�*ۢ�^C�,Pv�6Mv��ߠ��-+h�������.�3_#ιLǻP(�����5~��R��=�ͳ����}�#궠�&���]���W��w4R4�p�h?��ǳ�����b]f�uϓ���ɡ��+(ԗ��4��!�`u �4�Tt�% 8�G4�,dȾ'�kF>�!���M(>��/#�����U�#�vsQDN�G�t�7?�!H`�F�Iiê[��o��jTP���d15�U
�aWQ�~���e�(��VϨ���"�P�4z��������������X����>/=�� ��O�	��c�L/:9�C���M�<|*ڦ�F�az1�裀E�Zs���\<T\?�(�J#�)�!u�6�~ܚyHC�^��\3O���Cd��i�V�8�v����%����G9��g�cmmo��8u�"fh��muV��Y�N2�UO�(wT!���*���d�9��1��dde�U(��&����諠���/�����!�����	�(]�q�͠k��~/v��;�T|��bE��v(��d�)q�Y�L7�{��T����/٦p��.+�~x����]�z�&nܭ���W�g��LNE�)�[�<*A��c�(�X�y�S��1�~|�?����m��g^���[\G/�u�hڍH�����K*����~�!�h[�է�<�4���ߤUt�ը	7�*%�`WdC�P<�65��M�RX-c��O�#_�P�iHi�6V��<���.A���bT0y��`�	����|r�����4��\�Si'�{����RZ�烼3AF�d��1���j�Kh2��{��zA������	k$� �� ���dI]�*+QDPe�Y΃������F�*ڈp8br&2t�@�
ĩ%/���U�M�#@(�xD�!��"rɳ���`�:�^�q4uA��le�9��Y5
K�q��F4+Yo*���PD�V���_���6�1��p/��2&��h��9���EG1m3���!ٓ����=>���$��ob7�J�8�l~��1�M����6��?�U��_��3��lb���>�m���g�������ݭ�?�7G�Ӯ��������<�wc��S�Ǻ�c!� �w�,�l�q����0�Ɔp��ud2i�~Ô޽�el,�G����Ҫ9���'8�ٟE�gZ�)w���r����1l�~������IDB֖���߳�G��C'y�~�c���e�2����Y�F�l��ӯ��To���]�<	�Љ�����ͻ�ꍷ)�!L\y;4һ��&u-u�F�ZÙC��e5\(x�c�x8��w>ee�VӶG��LuQ#���kЙ���!�)d�jV��s��;�lՄ�2}L5�t4�])�U����?�Lh���������V�N�E��i����+�M}���߸�y�ۈ��Vf��o5�q�铚T.Ѣ>�h^R�&}u\�NzT���LU�C��|�94�C\o'��&lx��0U㟀��i�?Ԡv�G����hnn��9n���=��s8�~)-��h���T��f!�0p����3�13s߈�5O��=uZwu͌ �����]<��x����QQ|�`K�Ho�P�*���)��&,�-NV����0�>� M:ij��ّ�^�\�t�o������zE��y��+Ϝ���2����~��D4`)y5�/#b'�3�H����ĳ�:�Źy�<q���hڲt*+��p�E�e�%:)�c�\�"N��Ó�5��Y:or�y��N�6��9�3�YpI�Wz���5K�ڏ���"��W.����GF;C�u�V�5�R�f��vj��K�.��������a$&��dOf70�ݏ��H�p������#���h�ʸ�q(?��2�R�҆�V����=9qC{(�[4~
_Oo�Jv����nLL?�@j�D������R�]���\
�E�R�&�`����޽W�or}�SSOs��v(�=���wӫ;����Q����V,ay�Jt	�5�!��qh�� ���8(�����W��g>�9^�O�nbei��f�6��×��,Q�t����U�߽�rTТy��oauc�X�;5k6�L|�Z7_��vؙe):EP4�I�Q O�T�}��y��TUKE�ݧn0eEX���t؍7�0�$�'%%�|�2���{8�i��K�42[q���]����~偪�l�dr|��k�P������:=�uS�w�=4�,e����|���O�;���G��fQ���5���-�h�t;EM��K-���B��K4�;�V���*"T�᮸)����ȵ�]Z�$mnсNǩyt�'석����̨�}XCX��A�H�i|���;f�r4l���H󽚃{�W��{�s�r�A!����ޥ"�����!�����WZ�ll�q8�'+���3�uQi(m�/�@�Q
V��C��I.��E?>��Խ�|@���w9
�u�;@S�9cz�x�����u���#����K�)Y�����b�8��p=�Z��<���-Ɏ �>K@n�jȒ��N��^Ӳ�i��T������}��Y�Y����,��=�Ԛv����x�SVʲ�%��%U7�n�ɛ����Id���g�ǣ�|��A���|��MI9�^���t.��[�����7~��q��|x�N�:��JS�'�g����W��?6Z�}H�>lӨwus��׷�����x�N��8uB�&��&���?Q�L`co>���X����I/��q�{�����^��H}�m�&.���l��S�/��Q�(�n������:��~�ji�a�j��6W����W��v8׶�p��i������q�l��w��!Ƈ�ћ�`|2���1\��6��{��!������N� ��5T���/ϥxB�Պu���Ƭ���'`P�tS>w�P�6��uh�����Z�sw:�ǳ�q~���f�Z��r�5.�M�*s?%7ʦh�CL�!p�!t��Kՠ+:%�K�t�y|&�6��V5Y�xۦ�h$�
�᥼W��B��~��n5;��F�	�I@U���d_u������N�Μ�v�s�a}o00���2V�U�Xm��R�e�p���.'Y��X����v��+|�]BZǽ=Q���[���1�Wg��+h�+��(�f��G�Q�\$���طzĮ��Y��wM����R�����*�&H �Oݼ�߇�\]�7nݸN���ep������}�J�(Ζ��J�
�4=���D����{�;A6�<>6������\�H��� u̦Q�)��:vl]�mL�(��%���.4�ib�^���xۀz���}Q���A:..kb
�>u���66�?�A*9���z�}8u�eGv�V���#�=�l���.z�\)G"�o�1u�_��:�ċ�P�����+c^C6K#�uE��-u�Q���_�Go%�7�����_y�O_���}<{峸s�}
�3^]��*
U�>O�ڗ��[����_OL�{�Q������CP��|�^u�qN��!��p鋿ȇH�ȥ��It��S��G۫FP:�De�����@�e^���W��1������8{�O���C��y���md77�'�M�+�w<?�Wq����Y�^���?&����Xo���#��P��A��x�h#4��Zx\��U�<>miyO�h�l���Ƽ��%l���ZԪ��p�^z#CX���Fk�i�6z���Q!�)�]�	��JF��g��nG�9�H�X�M�S�[��ס^"x�����&�#��x�4BV���2N���CG锣F�Q�3�li�7�	��L���Z���Bͮ��s�n\����Q;���
�{�6�th0I�l�Z���0�Z���tF����{�(4QӤ*����K��%�^S.��-�l�81e�ᮞA���u�7=���5��>�d�ZD2�D̛�h��H�f-�(�ߥw)O�:��8�\���	S�^M=	�dw8�({�� �&*��6:�J��&L�7jY:yLM_���f�o"�8��M�ؤ���c�K�m�@��^�=./�X�[in�8A�����(����>a)Y�,i�5����l��Ǚ�|�>
P��Z<��)�"��%�lT�jsF�齢���K /��m{��W1H�\��A��"��L*e���g=��YӨ;=��)jq��3rU�E���Α~~���M78<br����Re���֌�M�[:Zu�D�Ǻ�E|ws?�s��&Z�<G�Xxp=�0zBa,��a��S46	,->�g{1��γ��:����k_����~�0@��������7�{��_������[x����s�p��i��a�ߺc��Ԅ$~� V��F����3/a��Ψh�j�	�L]����Ȗ����-ԋ���]8��s��p�b�4j	�~nk��<�.����H�#2G26O���}�M}=�P]" c� s�osKE��!�	#�35�����n�O	����8w�,>�w�g,��$П��?����A�F�|�E7����?����猀=�_EB!� �we�u�P	G͊��-�r�4�\�\1��@'�-�1<B]��5ŕ�%�m��fw+�홰Q���5�9�G`L��>]�h�fS�����8G>�,T�7���Kp(�W�q�@+�XFJΎ"o�*x���O�*3�|��H��V�IGT�c�FQA�k�`SMD�=�kO�Q2ŵT����6V���.;��Z�?W�CG)=t�V� �ӋY(Qg��m~�	��	^�t���|""�I$��E�
�s�t�>��#��Qs����U�����8�b�\C��JBS��֜�3�(�"�\�L_H��={KKK�͉~ܿ��ɓ���>$�e�?s� �f�
��|*#�&���3�q��)�`����^v�.��@f�<D�g��Q޳��k;���C���ߴ�w~/�195��F���QA�#���f�e5�P��y��8sv�v|����%4�g���k�0't���r�����o`�>6ivG|�����8�χ�x��D4
�M.'@���uULQ�8A!�(�F� ���f�*T�C0�`�˗$���Xv#�� O 9KУ:��<���8�ffQ��pj�_'S4�+<�B�5#͕�ئ��у��y���K�F�P46
�D�PY��قk�Q��+f�MTh�Ϟ��M���zv��z�+s�-�p��séT�-�(0��~Z�$�8����q��s@��@���w�cc~��m,?|D���s��(ڜ�g�}ż�O��cX����2��Ő�wa�`r =`]ѷ��A0���K�8~b��z�K�ӧ.�����S{�޷�Ѽ��r�F�T�.���	F��I���"�Ώ�����.�C?{���)EY����A�O�[&"�n��Ƞ��"���:uC��Z����)��������w���Y��x�(�:��N���tjN�bju��U;l�޸~�B��;��ul��A!o�F)�`��]��}u����M���u���1�yOJ�d��h!IC�ԧ�E�粡�b���5��6�݁�A&����F��J���nhVY`FiNEI�j$�|�r���gRN�Z���t-E�����F�����zRl��P���k���3I��ll����K�C|�ܟY����[�q�6z��v�m}<�DМ���SJ�(ʩ���r�Z{Eڂ��'9Ɍ����9�Vd~y�,��J� 9RP�cѶ�����>l_#ђ���~���=���6�<�\S�U SQk'���=9*���R�>[�)Y�g)��Lcr��z&ݿ�����2!�$�<���s�#��au}��$R	#*���!��_�y�~�UTy.������5�x5�'�F�/�������#N���SX�,ӑ[E8����-5F'��o��?��~���=|�g�LC3���⟰�����_���&�&��&N�:�w~�]ktp���L`��w����}�C�{Y�(7��J\��m:����>&���:�p��d	�w���4DMqڵQ�l���7�H%y�ȗ*;Ƈ��^bi��|�S��T�T��\����W�wWO���_��7hܺ���8��Ή���v�G���&�׷K[R&����[�06�Ͻ�C]#E��^+E���Ϛs,`�i'r��_$S��*�*�q;�1Z���-k��ЅRɃŹk$;q��fp��`���t�<i����>�}_�.�g�^W�f��E~���u�gWD���4�Vw���T��iy���v�Y��Q��� (w�:����C�E���	4������8��Fq|l� 杻P�=v�{'v�����8�+�L�
��ڹj�"�a���"O>w�"�t�d�^9@8�;��l��N�:cߟ99j�
*$_��ڶ�΍P���4�	T�?��dɢ�:kjLQDϙ#�o� ==Q������B.?u��v��<�k��11%���J���������K�ak�ж5O��[71<��s�Ch��:�����K�N'R���"��>.�䫔���0��ۓ��Y�����ַ1}��b�h���Nr�
�|���8r�\�O�*A��?0���(�I��}lp؞��h~�f^k�8lO��"�rMO�3�z��'�A�͊׈J�G�iM_�V����OO[�b�H��G�TB��o�E���\b��һ&Q�X�0�`(M��!kc��.R*����/�(��G��=����^خ�(W�ԕ3�>O`)z�U�@Q���B5l�?ɫN$MqQ��k4�Gy~�ëM�Զ��y�D��T���;�0�����q��m|��0�?�ӧOЫ�c������`76��Ҡ��T��Dy��R�D�[�W)�;������݋�1,Jz����s��6f�����|���x��@�!��<4AU�>O2ą�'�W*`f�.F�%�+�r���%�k�.&�f|Z.\��m||�B�.��;P�+��W���(�ōG���$�Qݘ�z�|�M�S��:8���e\���(n��=� �^v������X+5"� C,0� ��S��E�#�V�6r���)�ۊ��y]t�Z���&��y�G @ᚣ4��[nog���i��:�7�BWf��U]����X�]�O}��%��[7�a��y��������ւ���-'���/����:�_<��������e�k��Ŝb���.�S����1(:����Ӑ@���Q�%�g��| -�54h�ɡ�ۊ8 �N�@�j�>i���F�&ɚ�S�>S�:��B�I�v�il�H�v�0E�8��YD{�0���3W���e,l^E7Ac����
��a8/�M�J�XN���$��4���:�txk��8׹􉃠�u@`�ꄔ��VZ���-=��ى',��t��=<u�����8�#���*B-Y�C��{�>���eQD������v�G�(�O����z���U��"��S����ޢ��W�X�j���dV5UJ��CR_��눦#��m������J��;l�d�[sc{��j�r[ܧK6����Wl�Ң�B<�F�|��]|�����❫�_��o��3W�)����������o����|�/���������*��A�\�T�e:5��XXE2�FwW .OuWg��G�{ʸ�b��Q_���g������x��]}���Jث�|����~�DB����������	Q zSF����+(d�<a<����m�
j
I�Ċ>:��|_�韱���E��i$���?y��S�e�P�.?���u�e�;I��.�U��e���.�yP�Kӭh'"��ۡ��Wi:���mM�ހ!�(�hg"a��<���o��-*/�	[X��I�y�C�!���4C'Kr��Q�O���o�Y���s�EBt6Vi�����Dy�D� g�`r@�$�t�WA�p�}��5z=n�(=ݝ�[�b��K4�!��K���`K����4�m�Y*YgD�]�&"*٣�Vͷ2z��x���;#�|T�����٧���}�no�W^���AL���F�s��c�<���ŷ/{Ԝ9�4�xe���C���^		`�?;��S�I;c U~�z�S�F��@3����s��Ǐ���y���	��)�E���U�����̒���IgX �H@Tg4*���P�g�'E:����
Ԑ @�N��[�����¹�6*v{{�NU�r��5�x�9�ccc��t�[��?a��=	/.�?FY�QwIw�	�3���B��.���u?J�l�.Y�m��˫+����A�������XS�ק�����)�h;��Dz��c���;��v T��z�vj4�$Da���4P ӱ �r�@�c'M��N]���N#�D�;�с�n���T����k�EZ�8�T��
�04�ј1"jޫ����Di�Ym�8��&�Ԇ�E	"P�s#�6?1�{�q����EM1�F��@�-���kT�ce�{�m���s_�,�s��h �T�^uvݼ�ݵ���l�#��p���=��W�{ݸ��*�u��{YL��A�Jyc��A*�Z!���W�n'pl$Χ���N�D�?1q�
���*�Q����F�yf�vq�OE[wcp�<ҽ',�Q%8��[���'�]��F�@�ԂHiw7vLѥ�9C�e��$T c
�ͨJ	�Pu+j"C,O����N'��<�ͩ�5=�1�����?�	���C�����Jw:N�����2��Oj���<��M�P��>������+j��ca�F����k����|ps��)�Lr}�j^t����|�/�y�����`,3�E�W?��5���Y��"RM�AYv�:._�B� ���&�ө�°&��Q���ֽU���˓�W�(|��-�A�NYx��"�nٮ~/rsEg�v�7�4s*kt��lT;�w�>�>D�����p�m��N}�:��c'������W�|rO{i���2v�s_=z~����(�R���a��Z���H�"̒9���s���e0l�i�1"���8�Cy԰���d,�x�R\Gc��#�)��u�;]����l���=u�oE��p1�J9Ϫ{3���"5����u]=������h8P:���p6�hW��4~�� ���9=�������p�����X�Dno��_�S�#�X����ߗ�i���[0��Bӯ���%�|�Y��_����VV�������<Ɨ�ؠ�(g��Vz�O�E�`[����T6qy4��/�s�D��wV1{�	�}�K8w�2�>��#P�:߇��Mk���Fv{�:�c�q>�^��>!0��M'Y�z��i��<�u+�X[o����q��ul��x��q��\��*:�^��1����$y~W-#���+9�8{�3w�zô!~��[h4��G�4
����݃���n)ԥ�8,
Km1Sh��M�y��sx���!B!�'9���X�*���K�]��D9����#k��j��Y�("�7J �s��Uə�Φ�O����j[Yu�����D�^�㙕��L�����Z��u
kDk<r���,���hL)�l�^��8�6g�e�5��T|w�=B�[	����`zI㍆�Z��m�F���Qo4y�B� "Q�B2��-�>�T��-C�1�:*%_�뱑~k�K(P28���e���Տ��y-�B�W�MUܘԓ]�	�O���D��h=So���An����m:ea��k����"A� �ү��2���5	�A�� ���&Н'��bo�Pî��k]�N�y�)�7���1�:��i�6�pq>*}�Nj��1C�l�[�yҏ�>A���� �._���b:���}f�r���?uS�m��?Ϗ�L�M���RdX�bUz fE*�����1M&Ek���)O?^�B��K��lL��1v=4d����.b��p������5*�(E���g���xP���#8E����$�Y
JH\J�_�G�S�b����*��x��$�zG0�jݶA�L��l��?^�A�%���f��h�����F��}̬/�����M��U�͛`��
��뛿O�FdN����-d��{HF�?���m�|]�R��N�B��tX_:;F!X���c�ߋp%�x{��P��!d������616:�C@�ϗ�W��_�z&�}?���{4]x�+4�F��7<���z��q.\�D��ǝË��4�}���k7���`m}�
t_�\z���	n�����	�	��Na���Q��S'�9)_JEy������QrȠ����g�k�(KdX� ���dȨ\�J�E�c����
4�:y���E�T׳��f�݃�{F����_z
���M; �R��T�FG����Յ�~�2�~a��7wZ����7P�����KhP�]�[x�/O�`;�!ؓ���;`M��zl|��9*0/�w����C���sN:��(i����[U�<|�_c�DC������7[NC��n\�]��|
`�E�-# �+ޮ͙E�D�+F�q�Ds��Տ?������'�����6��]�%z�J�����E��M��Z�µ�~U�{�X[^q�SΜՋ��q���(�'J)'��60���jy���(�{��a����5��;l^9*3��Ӗx�r6�A��Xm�a�:��֘:���)C��E�-M��+�!@�ԓ�ߢ۱�(>SoW��?��[Q-�rr����N4�礒�.Jj_�x�����D"e�F˔a`p=]�}t�����~Ӳ'_9s���6�����D���-���O�tzz�2�F���1�?��7ћ�QI��Ϳ�?�翊����g�ۿ�kֈ����?���k�c�v��h�Vm�5�+Y���+�`�W5}4�|Ι[3��S���lb�5K]��j���`��(Vv�1�0o+�㸺�s%~V7o/b 9�ooR�v������B�����=$�26��R-���;\m�цm�o���yl���A�Uh�h4H�3�/�-�� � ��׿E�K��0�`�z�o�rܳ|�IP��:���	:��:set5J�&
��*⣞k�>7J�,���:�Γx��?���������o�z���o���nP��s��#R��	š��ٗ���Q�;�P���n�[�k��]�0����HMu�fs�6�T�@�y���V��tЀ۫��=����E���m��0�
���6
��ݍ��7�K�:�=.cjP�\)܉��VO����5#٧3��s%ט=E�US-�ԥ ��y6h�M�)��P��1�j�T�ذ&9�1�]O"����)��%kt���EѤ����D����,ӑ�>69f���	�G�&ժ6TH� ��Mk��so�����ō޳�F��LO;:ao� ������U$~��=e{��lԃ�ԥ�Ţ|�8!�7��oP���ɓ���Q��I��O��:<��n��-�	:�:�b� NOM��G���}|v��	<!_��MQa��̫c>�1�r���x(B��ik��eG5�@�'B_�x��h��G�v?2(t��f�T��E�P��T��f�]��#[��t���ra�6@|}m�J%`��=�'Le���_�y�5*˝\��lj�o�����\<ENq�Y���jv���.��h8W�d-��2M>jЌ�C�+�w�����sx����cp���%�.� ����'3���F�)������(���8���Sg/�h�����f�E �Z*��D��K>�ߋz�9��)E0�6q{aκܔ
�����Sm~�Ɠm��s'p�	�F�;�Wҝ6�8u�q0e���0c����:�d
�+ݝ�q)�+��!�ȋ	�����C���U��8���'~
�Q��Q'�����?JMH�eD�(`�T�<_}E��qv�Ohl
-�k�6��^]Y�t��[}�җ�\u����OR��Y9u�Q��{�ӵk?��P{TJi���k���j2E�2ا��ms|*�f�=��������K�0O"B�$����Ρ^�`������P�,B�+9|zzFt5<��94)�O~v&����� �A*	�j� �Mq�Ho��KH�m�H�&>�ω/����P�RZ�3/��Q{�|��w��k����>*�1lҳOУ�M�ܰ����C�(�C�e�Z���"�{�� S=�Q����h�,�LQiZ)igVx��G�౳��Sj�"}���h-�
��,l��f�Q@ң�Kʀ�!94.C��Z�#�A}��W�&�0��uϚ��T��|{�O9 z���s� τ=��s�\�k������N#Mss�L�Z46���T̸�r��ؘ���J�Z=K��1�J��dπu�W�l#� hN&ܸ��;t�i�ң6��7��J�xU�I"*(oӀ����gz�3pb*��>��S��ƕ�g>��V�gtw��*&��S��	B�4uN S�C(�]2NW��H׷�%���9�w�?F�'�'�kHi�F��W7�����J6���^,/b�7nQW(�M�C4�G�v@�����u^�ӣ���8t<��9=}q�]�OY��?�E���:�s��(a�j�)��`�C����<�O	݃=f#<C��{�d��'��	�����H�歫>ѺhiZUڨ�������:�7���7���>���_�gư���ѱi+������3�O�(�Z�y�s�-�fb�0��y�C�9�[)J�Y:��;(�Z���F��r`�rR�Q�����[tH��M�G_�C$X���uY�U�Mg4�+���Y���S��6�Z�q��ak���� C;Ԋ���.;L�j�X�JUzz3���8��N>��D�E���dk>�ʛ3��B�0*��3R�s�ҋ"u�΋��G��t¥WTC.�/u����������푾R�;ln����bv�BU�m�Fba���:���Jh6u<L�W� ��*��2"mq�*%߯�:�H�H�x!�{�xΝ�5J���y)��F���I�"p��5MjY��JG�Z|�?f��n�F��+sh4�NIZ8�:p�x��T���E�U'௺TQ�5�� � �q!�c>�<S5��F�]������&\i����wm�h��4"�\N�%n޼6�Jo��K/�w�����`ׯ��J~�I��"���E�1��P)ҫ�`���m��M��X(2���LTX��;?b��L����BW4@��ͣ�� ����Cvy#q��+�c*Ӣ���=���}�wV��� �4��~�Sk�F��C��RsD��?�,����gTh�w�w�I���o��9B,���^j;Y|�oP�����d"�|z�!�����y���4s�����[�[��mT�������'��6;6������l���e�۩��ŭ�U~��B����F$b#�^��;2>����qI��Lk)%�K/�h�C 47���qٚw�HJ	���Ζ
v��R F�KE��k�M��
[���Æy�J_�fn�@NuD6у���X)�0�x�`��G���-z����w��ϻ��4�@�D��b��
��x���������y36�z����E�����1{������SI�k;k���b_^.Ʊ�	Tr{V�W���~��V�J�	�W���b�#��*��
��{��td��5�T\�:�U��p=���-gj��K��uP�fB]�6*�Z��,���7��QY�}\[���b��b��Q}<}�v���-�1vl��s�h\,�s�V61�r�u՘C���y�_8ke�k�Vg%`h��+�I���p:*?���LQlu�Ҷ�nhE4�:��!Io(
��e�(e�U��m:OO&e`H�&��J�i�mޱ��@�>����hZ���[9�!͍~o܈%��A�7*Ba�C�V�Z�c�﬍F�qo�9���I2J�D� �OO�mx]��=^���Xyp��
W�g��?~�~�k_§�;�?���.#��"B���9MV�cn���f�7�]B����kzXXZ�b�M���g���f-b�����#g���/.cc��W_y/�;��E�]���0
tw��l��Ɂi��ani�>�
�E:9q�B9_���Jc^8هH�C@x�@/KCs����w�,�"���"R��O�q}����8Ȗ,�OR>�їKV��?�m�UM�4��L�|([�l���-m�h�-���e,�.�ױ�r�R�y�~\�����"����?�퍇�T
R�5KmZ>O��MOǲ�cu+������~�����Eܹ�!N�<�M�p�����b@jd���h�=<��Q"ș��sY����!���ƚ�,d�|��5�<�̳x��`z����$K�m{� *³��n��ݻk����+��Ve���ܟ@rh��U�//��D�@:���4�q�x�6v��+�<'a���ռir\M[���e�❷���N�.�7nև�gh#N���s=�2m�9C/�����-�H��j�KsV���;heTVѠ�TM �s�P�y�W �y��.Uj65��KK������+�Դ/e��~�­Ԫ���hY�E�r&�h�eE����戮fku�� ��j���4�=o,*/k�j��kgG��#�P)Sx�L l�2 ��I����`Oo��Lλ6�B�,�u�}�=r�e=�QY��u����2jj����vD���]n��͈҆6��p� V��}�*�p�n�C�}ht"�H,�����N��R4$�I�8�|N�=�MJp�zld\��yj��W��+TњD4�n�����Դ
��X�͡�Q�k��4���`�cE��m���5OF�,�Y�M�N��Ҳ���4�A�t8�L)�6�726nF6˃�['���<����Y�7�N!QD�lU�(�P�{�z@eF�{M����Z�����)u��s_��x6�h��s�O�z5���4^��6gq��ST(}XYj�#��{n��أ�)Sq�����.�F�cgӃw�*�Z�Z5G�h��� ӽ�Po��]�U�[>��)�Z��=�� a��Mk(�u�
F�X�)TDŉ��[�}�jLT&ek�g4��vT�%m�������M�+U5 jPh�`�g���#lu��Kuu��yg3�����G&���h�B�J� �A�;J6y��x}ۼ�->c�H�D[���_�����5c�CP7���y��ܢG(�7���P?�&\j6!��[�0@�Y��{����;�3P#P����D��ӗ��ET	d�� ���YTV^`���'��Y^*.M��|N�4n�,\_:�uz��K��^1�_�
���$F'����O���<X���j-�
\�iNO��np��TN�� �!E��9�F�Z�$��jߌb�C9]�h���K��	�y8��:E!�5AQ��Q�a���R����>�&�=GD�z@]�h:��%'ՙc�6�8���	w�^����ux?���mw>�;�}�����rQ���"�)^�`'��t�ĕy�N�����Fz����{�p����2i�_
�D��j����9�AktD�����9��q�x�8lX��_����J{�2ks�}����Ӱ���F����$���5@�m�#��G�����տ��3'Еә\��/�)�ǺS�JZz�)~�N���\�>ܞy#�)ӝj�s�Shq�N���)�SH�r�����NTI�2�q�U���w:9�ky��3˰i����lju'M��n�"��1�c�]�,�@��'�71�@*�`'�p�i��6�Y�?�`�u�[:�X�a���h�����~�e�'�����)�n�7��g��1�k7�t���SW(#}��u�a�T�4ֱVS-�2 N��qm}�����:N�}�t߭[�����^1*�z=j��ɓ>3�]5��޿���U��D����XY�w�O����?���4�j�D�{Y�x���oQ'�]y�y|L]��,=}I���+�kHē�P��Q�O�8ū��3�aͶWsU�VA�hu�"	�犖�PSP%����<�L[ٺC}��*34�<g.�簌ȉ��<*%�F���<b�G��u���`y�ʰ�>�8����r�����
��D���阍��E"�����m��W��h��5@\k�����>T��^�_E�ͱ��
�ʕW�7�Gܷ�F�M�/&
�E3a#N��R��Q��>]�S�%ǻA�jX�N��"�<s��r��Ps�QQYE��Ag�K�&/��߫ޜ{�y��vl���<������
�*=��֌��Ko{[�$qzV(T����m.o�����&nP!�;AϷV� =9�s�F�[�d#�ūn!a~aQ?a�����W��T�H���)MuZ*�B�#�R�B�*�o+��:��뻧Ae*-�mT�m����=ܹ��vۘ[���,�������z���̯����fH�߾�/��Wq�l����A6���и�6����Y:y
Mμ���Z�ݸ���6���'��m�/D�w�h^��A==T$>z��< �<Q��?�������8��n7r��T欉A %�5���
��5塚:BϬ��![�B�ʻ���Q��f���e�_ ��c�d+ا�QZ3�L}�	z�qjd�J?לt�C��ԉ}�}�I�X�~>j�Q�Vw8L��>)I0��}����c���ח1y�JĜ��࠽f�ɺ��r��lbf�&���Q��Lq
 
xP�|�=��x{1��N;�.<w��\[4��5�{���Ȝ����Pb�S����P��Q�/F����صP*��+i��'�G�i*E�u�-�xXo�F	��*�&Ÿ��i8�C�~Z=���F�+�(j��BMȡ�t!F�{ �j?�>�hz��d1:u�v���������ԅ(q�ݟL������Y�w�>���=�?ޢ�G?��S�i�p�e��	q��$efee��H���8�5z�4"Ku������]��IN����]ɸ�]�9�S���Mml]���}~{��"�*m�����Nu�U�BJX`��Is}�|)�-�i�7|��dr]���JZV�Z�o�/�G�1��������x0s�_��i���������f�B�d/:4ȡXڸ^/\��������d�GE"~���rM��?d�5�ks���\���2�N�#"����Ĥ�s_�E���!�zӨ��b|�8ғC�_z�@������Q/-�P6�V��B���c��
�<;�so$iz]����}���}�}���Y�� Hp�HP�,%�S~��`E8�6�p���l:Dɒ�HY�B$�M\��� 3=������ݵ�YYY��{�:�����A�D�;++����=��s����_�R�;*@��N [q
6���ۗ��ĬL�f%S�1s�7e_ª�Y��T�xb�h���[�������$W���v�l̘�4�bР��Mαe	���5�P]���:�__�|�=YB �
���z�\X]Ͷ�V��~A..�3L�`���?ß����Y���k��tC���|]�8����O(&��xF�+W �e~f^9������q?���\�JI�3���d��Ey�𡩭�@�ᓧr��%�UkfA~�o��<z��f�/�;� ��{8'�����Vǽ���[W��)˥��2\��!��	��6K0��R��Z��>��ԔL'&%{��5n���S[�Uw�z���F�lCM �fOT�U�4�������x0����~��%�E�J�Z��N_bc��k*�-�'rύ)#�NWUT���f��B���G5ibT�H��U8��͖9����K{��a�"���|䔻Cط1�A��s
��3�:�]�\�p+�k���/�������I��T�����C�Xi�<:��֬I��9�`ά�7�\��<�g|�
ڼ�?a�����z$��[�� ױ5�����?N�6m�r2p��s��-=<w/�%!]�?MPL�hhp�ﴗ]vW��r������9��$fOgұ5C�bA�H����K�Y� O�p:��j��%�M�����ZFf����VO�@�}������6<�!�-&����\@��P�s���r�U�t.�/t��$��511/֧E��:����/��Z��S�x���U�^�����6Ѥ��m�x��o�+�,�עT�̪���D2ꖽ��rny�*�HB���t}�yRB *.�G��V.6,ˁ��v��X/� �H)FМ�z��C1n���I�P�ͪ*:���^ 2  ��IDAT���lH�V�Mc�i3�m8��d���LR27<#�yc���8�d�QG2�=.�YUl:�����a���X2d�9��)0̧ɍm�CLc9>��_�s5;PM͸q�+#�N�T�y&�S0�|MEv���S��d>Y��b�
���lRJ���^{�����F#QI�fp�Z�5:0�N�|~iN�68�fV���]���G���o\������Ƥ>a ���4B�F3�r@#��qx�JЌ�i��F�F�v��Ұ�J�q l����i=�)���uB'fg�4� ���pQ7,�Tj>)���������ʒO�7�-σ��:�����lx��3i��!�=��#�f�&�р"��+�����ϝ���t�;����>�ֈ�4^W�L2_\{�,�ט_�����ԍ����i	���*�RKL�k T�@�)�~��	�~�[�Q�8':r��1���@Y~��AK��.�4�5w�$�yڽ2@�S�����o�L���+��Uy�g<�:��^-�>:5�_Z�$<�8�o�CP2��s�3)��\��N �C���L_�5�z�Q����
wU���jo.�G�{���cɵ�����Iy���3�Ҕ�*^�6a���0��[U8��JaP���˃�w�$����֞$g�jeff~J'$9�A�wY=*��N�R+-Q��m�!�,���qzOW��
[�u�t�2�r <x��S<ЮQ&"�qa��Ǎ���@�>���t�l^��)��:��6���ܵj_���S���T
m��~�%�P@.\p�J�~�c������iC����m�v*�S>+�B�0���n^}�u]����67�w���>��i-����������3)#���0�/�sIY�RZ��z��� 7�5��,J/W�QuC����C�E�Z���Uܫ�zf�C�|�����&����]�X���#y�s���r磻��*N*��Լ<v_Hl���$���� ��}�De4��R9�;�*�U�����U@����i7-c7�dϢϜ�=c��A6����2tX5���x�!�.Q���(H�[\�,�P�Ρ^+�!�1ö���n�G<A/�{�G�G{�򶍜?�Zw��kSqz��yN����d�>�� n�&�R+Ӣ�O�A�4�䜊��5']6��O@Q��i������O�6�������4������kqj����qi)�%l�ͥ�[�'�+>k�b���)4���n��ە[0�"��lڸ���4�z���||�n��lrF�vq1y9>�V9<i��G:���Jj.���.v�P���(8gx ����Ct(bQ�m8雒}��	���
9�Ef�3��Hj�z�֤P�:��65��+7.��ey&��ٹK���QGA緶�CvK���{���9��&.���`��H<e�����tJ@d" �`����y��1��x̲� �e�����ΰ�BN��$�V��L�g�a÷[r���qH�l�Y1-�6�t�M32Kœ*����T1���/l����jnBfF� 	���g��N}<�N��\��X53/4~t�4>�Qo�*3�B��;v�O;���2z:�d<b�,�9�X�9�Ν;
D&�j�9�A�B�>:0��5���ӎ�PȮ��tƂ:��KR��2=�d
(V�\Y<��Ryz�%f��;�R�����Ř���1W_��rUN�p�Ҁ�M��\\\��HP�X'�R[����w����OH��=
c#�h��e����j���I��ƈr�+!��b��;�",��e��G\�l`S�pۤT��ZTﲔ
�ۓ�O>���C&g.I���=ҖkWa�Ӛ�a���h�� ���d�~,�L�5?îo>GRt3o���ː�7�wvR�v�Od�5����Ɲ� )5j�]�-�l�2��hnJ��g�y�f�ٔ�1Kh�s�
`�łvs���fs�ȐB`�n�D�& ��S�0y�q�Ur9ɇםr�t�Y�i66u�8�y��u\�[:}����J]�N��Ca��?�9aI�f����Gr����w~�Ø��g�K��-U�ԋ���CY�}�*���W�����Z$@��ܓ�=���%�u�5�ʭ+b럗4l*�KWn����G[��( ����+/����{�;X�!�mJǍ&�x�Hn�|E�m�$w��k/]�ϫ
cӓZ���U���}�y����WJK*���Ĝ���8bA���L-�A�CI�0�����Ĝ���l������b��`���7[{p�!�ц΢%@gy� ��8����Q��9��c͜s��ю�� �~8Ȁv>���W]gv��{Ò<�?�`rZ^���5���`��65�"���?��{��L:, �W�5SMn�Zj���!���� ��T{$��.���.� ��K7��,˝?�Y2T����@��O}k���ԋ�H�$'5��F�6�)�˲��P~����,-��[���|����O|�� �8��,�&3�?Ź�%u~Y��nܺ �t��ȯO���ԗ�ťYoH�@�x���#�jMM��
�-˹��z�
�E[�55 �br���Ьb���(�j���njj9��̦�Em"�_��9b�G�&������=� ���^���j3uk�]Nz��F�Þv X�8�3�ۜ�h�p�A��JC{���j���I W��w�-r��1qI����ЫbO�T�v�M���)�����ن��o~��� |#��8�� ߁OJt*!Q�U�@�ל%Ϫ���@��>QB��{���HR� �/y��`��c���R�;���+Am���7O��Z���L"�'�)IrʢP����U��Z���QB�Z����:t�Rϫ��n��� $�� �k��03�$c[,]�)d��K� ����ɪ�}��,��	T��_��c"gYvз�;b86�IrJ����5�������}��q��|ｬ��ܺ�
3���#j��0�f�kK.��w�����8� �����^�%|����N.�M""��0��ؾ��=��FO�o���{SVS��_S~�w�N��>6�7$�(�j�Qi�!�lOg�;��20�A.nB
�F���G7����9�9���a�vnj�a4�a܉ɬ�G��1��k�A�9��>���u̙�l	y�U ��V�Ԑ��ȚYB�M�W^��X>�x��Df�/?I�%�Ic�����}�g6`�Z�V����/�.�_zU����r���{ߗ����õc	l��e
�`Я����q}��Wv?Q��4������^�$˳S!��^���Q�D��y	D�*���`�p~u�Dɏ��r^ ���0+j���ƣQ~\�f���y������c���s���n�Ĉu�Rn��y&�w�HNk.�r�Pꑽ�ci�Ma�>é�M�O��9ϓϋc$|ọ�#����&����P���ƌ�u;�d���g�^�i&C�;p�k�1�|>�D�Ȧ�$�;S0��s��H�:)�>Z{��>��)ϙ�ß���F8*�먶� ���,8��'9���*��1�|��:�W�,A)e<�_��>'i�l0�J�Ti��_���S�������+7��Ap��Jl��ݖ*�gz��I8U�fv��}�N%d��^C6�� $6$��9d�&�T<�Gݑ�וֹ˗�d��(� 8Z]�~3 ��d����t�R�/o~��l�K�ѕ��	mⰓ�@α'"��bt$�6���vG���xJ9��ο ��S2�2�%w��g��|��$��s���40��C��{ �}g�=#�S�x��e�w�ړb Ζ�����LH��F�	�8g����F�('���&�ڨ@ɞ @q�N�����w椇��������6J��/]������u�H�՗�Z� ��\�,`������F�aH6�Ѡ�Y�(������2��P�0#w��5�_���lZ�����[v���o�r��y�w����K<��1��q������+j�{�#���X=� �Q��S\.B. �Ͽ�2@!�M�L��u �|�L�.}��'P,�+*;Eˎd6(��`oY�!�z�ӻ��?�c*���H�#��i��T#3�*�c00��`�
!NS���؛�#�5�����}:?k����fpl�Dи7�ѫ�Ե9F�6�ev�;�~��2Ѐ��X���x4(�FE�h�@[Ϧ�qy�ܗ~Nr�3�i�}Ѩ����o�3bRi��nL�8 `�Q���8/��5�6ډ ���k��Iri�vS�\��e^�a�&�Rx�L�v�;N�z�b5�<'N5X���=��ciV�XvgR�$3�C�qvW�k6,�{��JT8�.34��4���'�M�ͭ�rV8���3�v+�1]���;@U�6�����8�[E5���:�Ȫe�~�����$�@�U�١괫�(t�n߭uv��;�ɪt��\p��97wY�8�H���4'}KF4����#"��pa:R�Z��˭,����x)���ΰng��nq�FV(���QQ/��q;�����!��"����2̕U9�ݤv�[@��m��|��-�i��',�N�3%��M���y�]?�mD�̤]�����s.gO2� �C��߿��ȧ�`װৱ	�X�Tş�s�I�ʖ9�����z<L7�H�f\��ǂ��1���᳡�>��C%G�����]��>�B!��;��*�L�;���U�ժ��*d1�I-�ݽmu��@D
�S�����(����7%���!�=ޔ>z_|z_�vk���=���Xr��gq���+�� �aHrr�sW�D� �s�y�H��r��8������|J�a�T�eqN`nnj"�Mu���M��N�JNa �q" �hu�/�O,�QK��2���0Il�CGx1r�AR��Ux��U��j�cِz����(q�TA<�����T	�'�]N�p�T*N��D�Q�C΃ٴ1���U6{�'�����||�\H���3OH𙏳ɜ��#�.�&3B~vWke�~'��D"���c4}*���w���lM�7���{�@��!�  �
����92�������h8�k�T���ʬf)2����`����9O���J9~�@��lNψ��p�;r���sH�z /\�J���7_�!I8*E�A�n˳�-�2��(��,��W���|�˸�6 �O��0�\-��/�{�%,깱�r{Un���3��p=C�G��{o�{�}��w[��� !��x��x���?��'$�9 ro ������VOeo�����(���O���ɕ�)Y?̪(~�Y���e�U&f��;� ���>']Q~
�{�����F���a�l^�J"׎J�J���L���p'g;�����I���ަ������K��{�༠R����� �<C`_��T���؉J;��7~� nv���-�ت��/\� @�ZR��֞��9m�if�����f<�ނA�XJe�H�ꎚL������f�4ú�ꗿ��n�`S:��k��������C�����/��Ů�����r��%9��um88���Z (�����yYЌ���pkOG�y�ɜ��DtB˳�#m�|��ll����W��h[3R�����٬�/�s�������<Y[�Q�lj6����2zG̡�	:��n�R7��p*mvO�W�3sJK�9�#u�V��Y�Ԭe���¬"��O��?o���o�^�ī�v�aVr���@v�Q��� �,Ӻ��Xvun���H��s�Ϝ8ov�S^����F�v+nMDq�!�W����?����2rh���L�;ل�5����4���C� ��乐���!U�0�WG#J_ѴG��= ]�����\���n����c����2I�$a�;ڰ ��J�B��]jd�K�H�5r�<�{� �p��C> ��(���%�sbSWu�6Di@�yR"�0��$�M��bl�h �x8}�󆆱��ء��'�&*W�G�|�b+���8?0/�S1D�-y����B	'S�y��6CL,x��V\�2-o�sWVsrz��F��|�=������@�;)�|K��|΃�M6cCffS�z/#�a*s��O���1'�����Ѷ��.H4�S��En��E������r���qA�4$5^9�?��?)��E?PR�ɱ(����ˎ�Y83�� 0�������6.�=:0�SJh0ǙF�]E�*�m�e��$(��p{z��ֹ��X��7Z:���j�T~5������=Z��H�$���+$4����X2ٞf��=x�E�\�pY��z{ʉ����zO!ZF4L`1s?�<�$j���;�iX3��Tr�I\3GK�1qZ�0<�@�<�ؕ���f!�]S𸁈���	��Ȍ�.9f����8e��th��t�}��͎>;�@;���#�����<�F�V-C��0踮6�C�f ��*H8N�`�S0�p� �nWO��8�G����)��N��5�q�����9���p_%�S����9������\q]0�h���׆f���|��T�Ϊk�Ϝ�����曛ۚ�#h���c�l���c�s<��hn�8�m�C�ԑ�SǱ�:����YB�Ϙ�d`Č%�ϛ����s4�����Ӈ�9����
Z��①fp����wWr�?�98/��+�z��W,ץ�ڧ��0dqyAV�]U�G4�P?��R
v�����u�w*�@v�8d/�e�sV7�Li&���Ӓn���YCVW��M�x�ܲ � �ˡk��Jİd�.�m+-X���=�;`�#�֞4�V�U:�K|���p������h��F���i0�����s������%Ϭ�ghj�U�n�L^���!��Zu)!��c�3�M�� �
�*<�h�*:�JR�o6t���+N[��7���֟�_����L�\Ŧj���U~u(��l����,;�}u�`Ă�j�t�["�8�S�i
FGi2N���(�ͱ~C�r���T������K�����3��8#��# Ίܼ�n~G��S�Q����tl贯x��� �ө�J��I��J*�#5��A��.8>;�kO��JڰG�e�
�5�	������ӵ�Ӫř5(�.0��p��p]�5��3ئ�ϒ�u�4�Xͬ�PA ?kh�26T���6y�A3�4S�P{	� �gh~�@ρѶ��$
:�)���fUs��1�������ڬN��C	ɞk0��-��	�vH���ݡ�M�$8ڸ��Ar6�{����4�u���� 0Ю�x��vS�A���Ya��@�HE��:���L2�L&�8젧v���U�a&_�߄�/΋��ݵ�w��C�>c����Y����A�W�I>{
#8�vK�Ql��'
��:U--˺qۼ0�a Ţj�����y�Òѡ�1��d7��O�����$P�KA��旉PX�p3wO4*t��fW+7'9Sp�4�Q��$�Z��	�Ԓ����Bd����@�޳5鴪z^��ɗ��5���R�$]8���G��/���`�Q�?$[��:���p�=� �oo�k��I��Q"�-�����9�j8?"v8顽>��a���^�N��'�Z��,I���}�TI'�9�;�z�&G�{ ��4��h�r0�hR��H��,�vG#?�!sES.�p��/���7�0�c�?K���oG`����t�t�|�%arqJE����0??���%5##�Q��E�XO�f�'A#�{V�+2T�N�` ��(��.���9�|�& �3y�)%F��Ep���L�X	 )@β��Ԓ� ��^���D��T�E@0�c�I}���?WrF�0�>� ��A[K�Dp����c�T�f8�^nܺ,g�3� 'G.�;`���%�Zd��A[倘Y��a�	�u:��=��s����Q�Ŕ `Ʌ���?��j��$�v�J�e`��K��əs�Ss�$�_��K�H���X����v�ݡ >l��K���X:#(z�䉮���i]'���Ϫ����jf���k�����<���#8d֖�R��-?�~6�	�I$&����҂�6y�sMq�έ��vG������	���h�"�����5�x��!ϊ��5̒$��k�������b�6��IM`wxp����㣜����|O Ͻ�u㐀�T6�#����+?�Uɯo���xw���*�'~奮=]��R>��In�]���d���I��f�fu�7
��d�Hy���}�cEu���`c� �:%^[N�q��]9�f�s�H��rs>)��Z:5�W��W&a�5N�B�C)��!��ch��\�: �n�W����⏆�5
ƩwHt�@p�6�q���x��y���k�`�3���Ki#��#�H�y��:�~<�ńOV��Ύ�`�K��$>�T���|@@X��D%s�yTWxQ+7C�k86��r��As�]����"6�=C3=l�cp�_��2�����Ykv`�)n���_�Y9�ےgO�h���¼��,�����X�,�>�D���O�	@A�R�Oa�nvv�4;�ҍ+z�^'���R)�`�:Z�`w]��C��ݽ}��e�0w֔t��9�����C��B*qD0��R^J%�r��o�l-TX p!t:L�d���#7��|J�(�0�k3��Xr�H���ٴ�n6��
���!�P���3��d���S���GF])�����<Ů{���mlPe�(1������23��/�h�2�;��ͼ�˹���e�/~؀�a:��6�0l}�9��`\)0��wqOX�Q�'iCf���T6�a���;.å�uo��Aۻ؋N�R���V2\`��~/�vk�u����<ʳ����z|a�3�ds?�ॲ���8��~���!7�����L(�O:�${�#�	���q�"$���c^8j���c��v5������3�(�@�(8ڊ]�.l���kUE�\"�LOܕđx�r�%�6帙���9|p���2�dI2�C9N��������E�>-�{�[�q绦����H��} �#D�G���L;�R��%�u��7���K0|]9;eD~ ��st����{:7��u;�����)'�g��9�O%��7_����7��GR����>/M,�����lP��w�c��S(`��+X�<S���|�ûpX� Ul8)�"�.i��Z-�h?����X:Ky4q��o�hB�H�H'���w:�q������%����;t>uW7?�S�������B$�PgO^`�??��Ό;>�ި6������r� y�&�,'�?]ȬK	τ�u��S�د�$�޿�\v���Q��a��c"�x8گ\ܓ���E��
���z�� ��H�a}�P�_<'ɀKfQ�X |��7 <�~y��-88Coܐz��R����-n7l�w8u�ʝ�'y����5�d0��&o�S�>����S%��ad굮����Ի^�7C�ڗ�m�*.�)���-98[���Y�`�8IkTK`�+A%��!��<J�xxx0*��G��V}�k��K&zn�����)_�{���:b���3���:F�/�?Ӆ̿��},��=���.C~?���3�Z��Z⋿;�>�3�
\G��Zz����gM����s����Oa���A����h���P�L�,��~ERsS *�ث5D��[�˚ �K� �#�U*��-�F�dD�g�>{(� ��G��ʞ�H۵I#���ήc�\�A뻁=�Ś>Ǧ���D�R��ݻ�di�"�_�.w�~*��]�a}V�<+x��v׬�?
���x�Z���"xk�a���K4aUnT���s��S�O�{zv���)A�����/��T+*�A�o:4�z�3�G�R�$�+�(4Nª���B���5b���hV�ݱ  L��b9]j����;*���E��)D. y�铢$f'���m X����j�Q[ϡ�z}-��-ʣ����D'�І��(�zD���P�;}S��� �$�R���r��W p�巾(�����c���ك�!����;}$�gR\v��C
�3�m|��
@f7����YMV��I�����@ȥ�ť9 �~~����Îs�����9��D�Br����<;?�{���Ԭ���*>M�:���ghc��ڱ��eV͚2h&i�L=U��r23�6��
��+��-���Hvn v6z1�g���O߷`��)Egg%ʃ '���H�˄�f˜��J�E�h�'�z�!݁Y
��;�ٸ�@0M��dv���R/����(޳j���'�HL3�*p�Z�x����9�0�Z�wI	!ˮ ��|B���/�B
��iqhsk���w�����}�o��!^��Sh�;`zC�8/'�!�^������c��XJ��Ff�WB:횴�iT�zB�؆�����|Vj�"�+�D���&����Q(�Tj�:bd\k��2�HvرJ:{�B�.J~0��7���,bΉ�4� �������l����y㭿.{ ��D�_�!8���@�!�ݗ��ܸy�fS7z�Y�����9Y^p�0rb���"	9��{/-o��26�!�O�#_Z�)��,	C&�0���I���o���lw��D�qj�S�n���r�d�L��m
N�X`�>^��X�����\�,�[RlZ�7A�3��̆p�$�9�\1�8��/��&S��G�ш���ۥ?�����<�	gM��=cfr��Z*+��`󟤏M�*8��x�$��z�Mu�\l`$��1y]U�g&�#����>} G|&�f�Ďh������v�b�u�����QK��D[I�7o�+�A��X'�p����?���9�B��H,q�Sث��N�T:h� #'ٚ���Cs����J��ΆTm%����~<e'*�-&����\����� ]�!M��R3f��10�)c�S���+��i�� :q/9�AрagNWl �Y	M����z�>�#��|��dRKzl�b˝�)�?�q�@P0n"R�m����-��!�N"a{�%:R�}�l�0��b �V]W���H0�D5��3smr�Ҩ	�s!雍!�&��H��O(a�� ��-|oLZ��s��z�Xc�=���MK��Sxz9ÛǮ�+�3��n�׍�����Y��D��'������2������a��� ���d�1��"��*́D/ue6>g��yG�с�R��Tp���eqnB��n��..[\�FC:�"��-]J4�{Pשv5��4�2���GX��$��@ʅ2�O�?H�P��L^R�Tp@`��`���v����V����Z�h|���i���5z:_>[�+2�b�r,S���6�4KG�G@f�
�����P
���G#I�RCż�g� 4�:ή��φ�(�2hw�{|T�5B�O �&ֻ����0\��*% Nv�ӆ�2�P�}x�-��z��W)�$:m�=��=)��RR;�+5N~��^d��1�.��qk1�q���C��lt��a�T��$��ZF:}�"�ӏ�����[o�;�O)u�K_xK�'��s�/����k�īo��~m��f��<��WVe�H88)G{Y\T����`�}�%�ݧ�_3�	-�����K42Ŝq�^��2l/ŗ�y�NV�HG1~� ��J���_�DPL+��*!�&
������{�>xǜBۨw\:6?kh����	&�����Yv�RΆ�Dx�Y�&������*��Τ���)�2��þe`c�����P��l��(�g�A*塔#H96����~�9�YK�X�w���ņ`�]gàO�lv�~������|�1����W��'e�T!����D o �5%
��1����V��yn�݁�%} S�+�Z�y��_���<����A��ak㢌֐
�Nm-��)7_X��Gi��R�BE�<�D���k�S���Tʮ�Ǣ>���ѧ%�H�O8���|�VE@��\7<,m<�>}��V~�.".*:bF2X�J�v{Lg�C~ l�fDV.^�1���6'fbʛ���rѥϽc\�qH�^��њ�[I6e`z�i0������ߖ�tN�S�P�oK�x�V8���99;y$7/MJ
�\���+/]}U⡘��9��N5_�X ��H�)N�ga�l�����^!��/l�V� QG��\�òC��nH 6'3sR̛����H���"�#5y�t��b:��,Z����J��\XDv���_�B������'4"<9q���Z���	��S#�Jo�i80��.8u����)Ĭ'��CQy'��8'~��h��)%�GE6�=����(��Ԧl+��M\�a�zF���pL��S� @���Rj�q�Q�����c���k�ڿ��4`l��))d�r��y��t<Y,���'������mk�͜lf۵�:7y�0��1�������������ci3�����7���u�䷖�==�b�*���F���"~�/OnI�U@F;44{CaZc���3�ǝ
�x�w����4��F����
�(5��C�;c��ƥ9y��<�7����
�*��2D�=����j*h��8F���/^�2�rG�U3�:T�8�g������t
�hz�X��y�{�V^�ǿsMs��st�:��<���	��e��Ĉ�r^- ��©v��lx{����N@�7����!l`Y������I�4�e5�R�t�*-�t��ao ���I���V�*!���&�-ϛ��3�j��g�'v�fk9)�g�2��{��-��<|�	�N�|Ws��(�1%yȑS��0��Og��%h�53���j[|��z�>�:�əYYY����i��,�~������.�f*)�_}K���Oeo7-�ȉvچ�CnÙ2{H��|8�l6�5Eγ��u �?w^V�N��,�	�.�t�<K
Ż���Ƽr��%�1l��J�1����>��>��Ҍ+�x�aT���*I��]n�)�F�n�S�T����a��OiO����wJ�7�#$5���s�;���m�����p���{��� �[����$J��e��Q���� �K�bŹ�H����"S �Y�3�qm���j?)$�����WK�����������Uf�dDڕ�&��򺗗a�gqy�K	� :9%�v��tyq�6�W�E�N�V��������>����^��s��LOQ]B�m0�*�Z��귒'h5�5�e��S���	�v����k�Π�:'��b(mU+��&�ML�W���A`VC�f8YvD��#�;h8��Xp3W�dU
3�ݩ�Þ�8�ک�agt�n��5,:���ߡ��?ó�hײ�-v���ڹ��F�&R HbK��%��P��T���/�6vk�۲�z]��洴�æ�8���a��{����,��m�!_�6�-�Φ�X�,̎N�e("���r��d`�*v,zŴa�8T�p`�4�:F-��	Z�@�0a�G�q�<�~!�S5����P$�M(�@����6��l�PI����vs�6����CK$=���5����G�帘�ɉ��E�0�`D�J�����ڒ?J+?�����"�,#�X�ξ8C.Y�w�{��~�'"'Χs*�)��^��v���T�7,~l�8���� �Œ�������Qܧ��'p�ۀ�fC�X��o����k�$�ħp ��hEtA�Ĭ��l{�����\Q�s�a:S�ATn�ߜ�hfZ��y�g�R��(P��5u�,�x���sN�	�|*Z�1��U� ���, ȡN5�w�ӎ����2a!w*	>�gV���-Ցb����c˃���E��-��ө�x�~���}�,2!�	"B,i�"�2\��z N0��Y��p�Y���uqA._��~��OwN��{rxp,K <�4ǯ54K�hx�L'�[4�����:Eí�=�0�������R5JЦ�~��s�$�9�g���$[�ɓ=�8?�=${��ڑ>�A��P��Q:��Y�T��l("�όώ�<�U7n�Љ#��L> _�\g\'�;y�5��1�K�
�-���ŋ*���s����=�R�����cv�r���i�T�SI���Uz�Ef����������8AJ"qݲ�];����7#uv%�
a�Sӓ��c��kn�sʟl|�,����{�R��ó�=_�O����&�Ǉ���û{�J��14;E�֡�9��t TyN*��t
ǅK7�h�X�<j���y��@@ع;�юF��6M��@|��H�*m8�l�"uKG��	�Ɨ*E��-���1"��w���I���_��� ��x>m�:%/8Ɠ kw����B0�;C�\�5;P�SܛY<�+7g�^�� j^ Fa��;����,���W^���s��rYp�щ�$'��Ǹ�Q�[*4�F�J��Z*�8���eq�����y�}�?R��Ѐ�"��K���Q� ���I�;-U[R땥֮��r[+�@�����<�4�0�Ǔ�H�j�K��3�;��dcs]3���ܣ�ba?lב��/��|�oi�[��_|��*8>3=���|�7d*��*�P]oE��JҐ�,��e����bv]^�~���1��p)��<�#��P����?�,�?��7-`?���q_�O�/���$
�+��� ��Pl_l���X�2��\�b	 �8�V���g�sZ�}+lL@�j���1��8�C�a��7L,�FC���@�x����a3X0�����2ć�}g�C��w�݈��ح�9��?��ʋ�}�_1,M�<��T�����l�:���^��lk�Ԋ��A���3"������P�\�J������X[~�5�'��X,��?8;>}��m.EB^+3z.o~��N��<��vG�^���6�������N�xj��W#�v���[������9�;�s�+w�Z�Vb��_s{¿��4�p�m,��m8l�<ag�3������2��o��sD"7(�~}fPh�~�I�J�4�
I��7
�0���,.]����H��-�bEu���A��8͆�U,Č^K��	��Oa����k��&:8^��T�F�ɗ��(�T�H�CZv�����F��H����{��{٬�ʵ���@�o���k�"��|��S�Tq	�,�$�rvx ��G5�����!{�MY����Z0�nѝWBp6�aNӡ�#�*G�%egO��	"OBH��2�u9+�0���K$�\�Ԍ�p�e|OB��O=�s󓒚�Ӊ	�᏿)���8��veB�{t�=�S��S�%u�U��V�"�z_�U��UQ�h�7����oܽ��73�n4�l<!��`�2c�h�gv�R��2�D#<?;����N�GXg�oNL����ÎK1K/$=sb34,�p �)��I*�)�!���-�t';���= ����I�K�o���9$G�`W���@��pN��XёYG' 2+�w@��c���J��'�m�emk�">f&�|/�.����HM���}��?Љ38�&#Jm�p�6-]t���[�Ƹ͒���zS��l%#�UU8#X����cƑ��J4ff�iʸt�=��M	ERR/�$�K���* ����}�(��C�c6�,--�3#�! ��0�	�s~!A_:�}�T��w���3��|`���8G@�Ϟ$�NO�7��58�yuT�%b)���躙u�301��.���1�	.��ⱈ\�%�MrN�YՖ��g�x}�&���+���)!�N^'��|]ܗq��8��OY���+��{ʁ�����hɍ�^{�Df�������K1�xn���"�O���_���eyج �LI�\3���9;�!P�˃{����$��=M����a/�
p�N�a7�K6�*���<~���;�Q�9h5�E
��*U�]eKzC+�HB N �+ZN�YN�ze�p{�H7��Բ�4����|�_����o|�$�} �n����l�d�L'gd.����H�ik�#�ҁLǂ��h1d��ce�%q}I ��W�!�6�fR����>+f��_��������t���[z}��I�񬍎�=f�K>9�?�HwDI����8�r�%�kv��4��<^>˔p�)�ߑ�̱<y�`.��䖱6����p�5�H�=�!PY�����MV�T��=)R,T�T9�G��{��	>wN��_���1���k��kyy��wenvJ���_�yM��T�UKP�߃�d3	C�����i�dRVE�WV�˽�Grx����U-UfN�`�Zⷪ�M���cpH:yW6�C9��{����W�:���l�����2�Q�I6�i9j���:��ϗ���g����?5��Ɇ��Zqﯴ;��ܞĊ��"v���pE�m<��+�0Z�7��V��%��;�N���s��Гx/Y�U�?�i��~�Q-�t���j�R8���O����W�ŻYwZ���N���a��zC�6����*���^��]~�� xv�`gS3�Ͷ�O0��{n32efS��_�}̝aX-�2v5�rXM���2EK� @`�y(S�ؼm��a��erʥ�:X���W������ "��KMF$�Io$˒0'q�]6���4l��/,�L��P� �*�O���nl�`���C��`ਥN�
Cˍ���+/����w����-D��S�:��Uk�rjN�
,�F�ZW����'��N���ua����,U�uܲ�ہ!J�3!'ٞ�q���� 
��<�R#�ȋH�"�7e*� `�&�_QN���Y]\����ev��UDq*����������4ke�hM�i���w���q�h\�D���#�ƍ#4�r��t�4zZ�$�c`6������' ����]���x�(<���2��n�F��-H ��m0Z</��f2z���g��] P7o�$�hH��wT7-/��܃�>�B�-����p�-�\�tU^�a�>Hźjq����udn�`��(�Y:ek�D�p�q6;�	,NMȹ��ri��{��GrR����r ��3�g xK�j��r��:n�>{_eX� �i4�

�8=%��ˤ3�I��GV�y?ŤD�1�yQ<Ն�\m`�DBXS���	�R�8�tXܞ��3��w;<R�0�8�	8�B�L��H���jܐ�ݘD��,y��Rs\f��䣏>ҿ���+ڠa�n�9'�>�^rg�f��Ӯ@Y��X�f�� �e�qZ9m8��Lb������xQ'��t&����f�Ln�C3�\#�� ����]r"�?w3����e� �p/fR)�'gg9,ioD�~�5I,�C�[���˓��raeU��LϜ���^Q=��>��4�%��	c�X�2���l���bL*ـ�,x8O<������V�H���N9�:I&�|�Ai���wEB>��F���Օj�"��æj6>�Wfg�K�w-+>����3������}_�s��O�= �("X����-�u�r��̈́`��ac�S瓩ĜL%�VhK��p�p��,P��d��'�lk �B�e�N;�/�A�M��6�qM��޽sWl,i&�+E Ȏ�o�ڰ���tڬ��`wG����?z�N�_��<��9���b�t*Ǯ�{�z�}J� �2\��E��l��DL��3<��+�yS����Y�lZ����,m?A౱�-��ΩB3]�
J��T)�F����ή�<�T=�B��uK�)|�:3�q��Y���y�����?�g�.o�|Y�ܐ��ɍK+rneA���}��+ҵ5e+�)-����^���}�F8�.�{i<e�v���w���7�����='綨b�TRT���F��ڐ�6$)0� �\k���>�Xf�B���5*A�?�tkƓon��@�?����T���	\q?��w���o,���\+\B�ߞ����-�s���Vqg�^���J�俇�Y�'S����������
B�� b�n�Z�=�kv�����|���-<��;�/]H���8����:������3�k��ͻ������W���o-����7��u���w���>;(v,&Gt��ȘYr58ۖ]�N�S�v�T�)n�4�1t(����)�?�q���m��?T�q��7��r���*Vm� `d�se�*�l�x4W�T��
gY�:���q���+rZ����3D����v>�ezYT�f_�� ��	���;+/^�'�Z�#91)ǁ]�8�N��#�VY��@�bB��%�Kʫo���R��vt�C�ݸ���.e8�N��݉$}sHx��Q��/��/���K�޻�e�1)�~aQȟ8��E���~���>�#�%e��m�";�6?��c�����H)��A��c�ȩ1F�tfH�1�?�h�����(w�1dv���4������#X�{�w��X'z;�,#,8&�F�%m_K�<[�Wȗ���k�>�(#a�������T\��@�Ee^ n�����LOL����Ir���{%q�|m�|�D2/@���Բvk�<C����&A8 �g�7?����ܸ�zaSgWku9L��8[7��㖅٤N2�d	�>S,J���H���˫X�	��wc 5�VufP�JX&`7�N��>�c��o�c�3j"��:���N��Q�����X�T�ߠ�O��SبS:+J��W�_�o�3*ٳ�|�s�g��_�>�C��dM��
���T�q#�3A٘'H'S��L��@@?��1%Zl��`�纃c� O����c���_�~E3kj��=��zf�.` ��U3��H@v2s�1�K�#˾�b��5y><o�_�	J�s0�Q�1_���3z~�9���М�S�7�xC3�̌�;Tqr�p����q.�dBn���
�;�.|��KxƆ��VuG�?q"��\�:"K���*gXk�<��K<�'�FOr ��|E��&�����$n�� 9�Ju��R��Ԋ{R�T��2��]v�7�֭�r����=��5ʅ�)�� 0z��q̳�ܿ_.���k��i:����� ��0�ϔ���z���EU
��(��a���6l1��|Q��g2Oi�Q*�$�������,l�J�.~ ww�"�9-���dOܰ�g�i���e�x�@��!�p��g�DG{�T���n��=ۓPث�<א�k�]��f+|�Rw�c�\X;|��J��C�P��	�'�:D�B.+����3]ϔ�a&�k�գ���H�ӬzpOp/�N3r��}]� *GR��p?f�)�8]T��J} �<��l]���kRĳlVp}^��m�K�VMnf�Pf�5A���.����񑆑����=�A^�S%�H	H&lZ=�2�
�½h�~#݃f�խ�ԍ?(z�f��	�&�S�/���,��]���8��=�-�g2G��i��^}0��w*���8�'���mB�<���������F�յ�׽��(������;�	!��ø�~!�3|��b�_]�����,}��a''w:��o��g�����H>����/{����&+r�,~�=���f�Ϸ��7�/���>�N�KcaV��Xsd��"�, �^� �ڭ҈�c���6��VM����
9�/b��P^��9�vvB������%����
~���ؠ����4,% b��g����>�B�HB0R�rk`c$���3U.\�&��o�kD��er*.���Yu�����%�~�%�ZyU��
�wp�z���r�K��ѯ	Iw�mH� �N.�!9"1���b�r���r啟 �;�<�L���`X�K$Ly�d[��x9C���7dn�2���B:��{T�Y��� �J�U��z253����S��ՙ�Q�Ǔ�ԈO$4Pj��,LF#H�F���#ܱN�I�n�!4%eL�>uߘգ�d�������a�����;8u������ͦ�D�������8�.�ć�?77;*g�C�0G\�:��6tP���Ւ��%ټ�^q�\���Ta�7�ݩ�˯|E�\�.��:�dOz�8W���<�r|«\�rvVʙuYY����8Ϟd
5�J�\>?'q�v�,�Uҕ�� |����������`�����f�}~�6I�ݻvrz,�v���� GU��D�@GD��:N����ԅ��4E���F�?��p��x�N_3 5	h)-4w �#�W"p0=i3�IJ�����4{�\4���@/�7������#h
�C��o&��R0���������|>��͛�4�~$��:dy�ԡ$%`L?I��r��޽�ұrm&�q]�&x-���TjB�
�V]N���7�(Ϟ=�5e���)��5L��������/�{��1K
���-e�KyUP�5����w���a�E�y��_̮�9j�ݵ�Ni{l�[��8rf�>��}�ѯ�	{ғ�iM�_��Y�ܺ��Y9�ّpV%wx,{�{ =�څh��d}��q�y��vI�-ܿy���������
V�������K a��f�hueZf� 6��-��!��	�r�	�{�u�~7Gs��U��H�af~aa	 դ�4Cq�����ܒl�P槔�C�hJntkIE��=PM��/�(���gp��N��gR(��%D`�`��L��	"ت�k�;��Y����U��g�>8T��kW�J��f�m�����j	>���l�`�̱c�#`�w:���t�� �u��g�۔n{ O=�zK�u����!f�����ݏ>�f�[{A�|����� �G������n��e�eչ$�d�&�^n�������׮���vkk��'_�ҏ���zW���;JL ��^4ac�ℏ��������[o�!�~L$�v��,�L=����W����f�j�ٸ�y���q|�ņ�d���O9����h䨃]�{�]�[FU5�9��>s���w��?����z~��=�S����}�,y<�buD�?�\9�~���՟1,�c�-��bY�3#���[}�s�*g�D޷LN6��gR����������z��ܵ�C���L"Q�Z�m�o"����2y��R��_����8�r��s��C�(�@2Pbp���,��$�66���ݠ8�h*
`�8�_��a��G��3H�,�;齷���j3��=�3��ww��+,$0H	�RR�$��~��"H�� ����Y;;޴��嫲*3�*���sov#�FH�49Q�5UY�_��{�u�Hcq�ѡC�����!���t"�dP�)�7�����!n*#��$'q �O�j�����SD�9mb�Q����Ϳ������XWmA!�-�Ә[<��(�D�(zM)�u���M����(�B6�ǟ}N��:|�!�c��$�ν�>�t
�.>��3�xH��YhЭ~�D'�0���RwHoH�0���\���d������{�l�JN3e�W�� ����򸰟\��m`X���\�LTy��K�6W�`wg���R>@��%#(�_��<Rp�숬��^�d� 
7���W(�������(Q����{�xG�,�\�N��L�ꅅ9��AAu8}�gN�O��{��{��J����]g~�pf���E��>"�N�/�������q�6��8�/L`�ʠ���"� ��|�������O����l�p��a�N.>>��w��^9�k+���p��]d�Up{�I���SϠ��aI&js����ΠP���Az�m�8d^��X�&cu��gx8�1 Y���.ޛ�`9�Sk�]~ �~�f�ވ�b��8m���d #�}�AЦ�qK�pp�T2q�����w`���[�+�����A�2��/J����_�O�!��8!y�ܗAy��"��f�rPʵ
@�9����g��Bv	���������Ke:ŔN�^�pA'd��T���R{I�ʤ����� ��eqβ�d���eo���3�
 ��+Y)	x�z$�� �D�X��'	J�Gv,ut}D�Q>w��\Za�1bs�~��XMm�==�S'��n�p�sh���a0�NO]3�Aq_'[˥,���γmVj��*�$���GQ�7�Jp��4��.x��3n���5	]��{5\�M�Vtz;�T�Hl.}��(L�VԶ�W$��LB�<9a�i�}!J8��>��F�<ĳ��}l��	W!��S��=�4�E	vl�x�Cp���x��Wi��x��al���=} �w�泎���'o�%0�!:�D�p��a<���P�������X�N�u��dj=(r��
U���.Ap��+�p>w������!�F��������(�,�x�}�U�������.�>?6�[x��W'��bZy�gu:T�~uu��YҠ�������T��VF����=�RE�0>=�Ӧ�]|������_�Yt���wn��KV��s�k�J"/�r�I�4z�{��1Ѥ��-�����6��(׮P��\��Q�=��;�n��0��s�A�^ G*ɂ~O���<=��>A1�B�=?;[�M&_�������Y������lgu��������]�z2����N�o����_vG���s�c����3��w���D�έm�����-����9���>gv������� ��S��+��}�/��Z��h���z�< ���T�Qoh��H*�i*ښ�̂��@T�2�t�����C*��L�FK8ä�TWMBC�/����R����4Z�L.��2Tb��jͺC�H-�b��!2�9�q�v-8MX��^'N<ʯǸs$)��C�ׄ�{�����yp�������-=X���9v�Q�4J��B{�$#sF,I��w������F9�jj�N3&��f72I�{���3�ܤ!OW�켶v���ʠ~��� 6WW0S \ꕑN�E%�ȳզ�L��6�Pw��F
6��_K�F����.�uP3#������OP��_�8�C!��LD
���ת��砏l0t"d�G Fzp�����Ϋ�=��޹H(�ݽ5��-�[��̋*Xt�����9���d��[.�xOX���Ⱥ���(�	�no��5�a�vy�������r�N£`!W<$@�������'��U|���}��n�`�5q��*� xc�]���VCf?�ٙ��ǯ�%����\B�"{��Gjg[�C�GS� B]a0?$A��OPL�.���G
~�Gx��,S�"��p�Y(�!�n�rg��Վ���-��	d:VD��l���k��F�r�É8�r���ZJ�d$%s������l�\�ܷ#���G��P(�݌�'�z3�y�p���T*hVX�#�B����w�����0h��� ?��}	�������n_܎�@��C��&��:D�V�]򽔄�|'�IZJ��M��hFGJ���+dy]ڟ(��h�J����^�Z�g�x�ל�(oĶ�y�y����������k��O~�#�<sw	���Q# l����/ai:߄SN?�yX
{8�3�/gA5�"�i�>�ǆ1�=���Q*�0v"���E��N{�,..�m����#4��k=q��~v�\�|�sGp�)�
"i6��Hހ���
�A��������ڬ4������h���3��`%�4604������$�{	�X�y&�U��"Xw��(ePͤ0�6� �N��Mf1�"s@�E�(��6�_�0�c�������+/�vqlq�6kQ�1�d반�mV�p�Ƈtn1����p�~���W�^o���&�"X���&
�oW�e~>Юԫ��x(p����p"
7��+����ܧYL1АJV�)�<��,���	rOʹ�-49r�ô���]��!��*�E}��.N��Gi�������/�Ԓ���*V6��G����������w,�M _N��3�,���mޓ �����C�?J�' 6�{����s��O?���;[���ɽ����1�]Nk�Rn��=����E �d45ڭ����t��nuqa�n:��;���g���u�G���{���_=gz������K##sͿ�9��
m�w��֬��_������?����P�߰����z����jI�/}�2��$�F��%�h���&b�"d��D��fB�Rj���	y��Ёz].�������# y����v��B0�P�4�+��LC��D@�Iy����hw�4�a��[���'Qn�̓è�eC�@�Ag01>K�jE��g���V�*,v:0���G�r���t܍�6�ױw�>Jwb,J�=�c5]D�L �H�e�⠸��������2"<93���e�C
�=
�<4a� 2�
��6�Ms�oU�ѴV �v5EP@@�跰��7���M:�,��i���
�6�5���AZ���!j��:H႓����H/A������x��L�d�ϫ����4��nR
�'�B5"NX���T�:�{���ئ��A?�`8E �ds�nF����JVH�d���l�%��������UB���XY���Jp�CRJP�s���
%CIe+��2�!�z��J9#�������w��3�����B�N���L(|~��hkɕ��{xqza�?'�Q��+�_U��:�Pl4�D� �{x��ϲ��kZ�j4Eެ��f�(&.�`Ȥ+�ߖ�t�rX� Q(0u��B��٬�ƞ[�PsY�^:�2����G�?C�[ߣj.Қaw�~�j������.�UA��<�:���Z����3(�ti�Hi��&`O��d%÷xl�a�CKur�%�8�GYG�:���;�WTA{�T�hfE�X,��l�Q[��NC�=�V�^�ADJ�>d�u������$�d�u��@�|"�'�7�����1�&{!\�~M�;��d_K���F߻wG):t�+��B�JE�8�}!�2�@2q�ǁ�����3I{�!8lbzBȅ�=�/\�TEv��/8�'��(b�1\�����`3�sb���p�19��V�À8@@��u����%[��~h�E�������K�pnn��-������$�������Z)��?�|�hKpx��9����������s#��h�i��ޅM��G^�<_��Î���{c��n��Ď�7� @Z���A,�A:y���	����
m�I/l>���tr��,�1�������z�k�{X�gJ�l ����1�b��K(2kc_+^�9�wRn���ͪ��"e�S3�ٔ�44B=�{�`)�u'ϟ��x��(�5K(*"�֯)[�'���p0�l�tQI�����v��m�O���_{�U-Y�>uJ(ig� i��ą�6�E$&vE��$ȯuF1�=��� �ĂJ\�t��f"u�����2�mX�]�̀Ug�5�����T�����[{��g/��j04�6�O>�s_L���u��|����f4�x�-Sɮħ<K���A����@>��<,����17������R��y��=�'(t�Ԍ���谧=>���5�H8UwФ�N�`(4ӽ0�[�.d�i>:(�j��*Uh`"PS'�#P�]��|�H��M4�F0`Q"by�0��I
{�Q��-]F�J)�u;�=/ϼ���	-�I_ZV<4a_�K� �
M���T��E�q)�A��]D��a�$y}Vy�{�tV4�l��D՜������3  �dz}4h�ܪ���2M��;/a9�"�5!���%[������=�9�W0��tlJ��hP%u�4�.���g��L:�-�]IC��>4����k�\7���T�$��~}�r�X�6L���Wh��T����ZG��T���fd��-�9�i7�j�i��x�D3��{�k�S2F����N�P�DΏq��.�ɉiUk�i]��Y&)�>2dd�{�$��j%�6����D����,���\�.�v����(����K��V���4��8u|A'Y(���Əc<H0��J���.�Ŭ*��"y�XZ�F1�UPt��2|�r�G��e�F�\��G�������1���اϗyC:u��~j7k
-B�^o!�)	r�[��^��@��dכ:�z�w�P㿁�8\�	����������T��J2��=��{���l��l�w`bb
{��N������t��s���PY���v������>|�|�	k�ľ���*#�N�?q�J�{D�{�V�t�EǊ;fߔ�f���`(�X�)xT��hX	�e�$�=ԉ��Ȱ�e�D�W2���X�we
YD�,Vx����hD��$H�3?��^Q0*Z�%"�)Ŕ<��\x2�Eba-�CPɪ�-�3��된��1���*�V�u��t����#�	��[���a9��m_Q��]�̽F��7��m$�Cx��"�ݾ����������3�tk6HH��:N�p�o��v�O�8{�4&f'U~��;N�� ��&gG��IDLa��"�8T.�I���Cu���1�'ڴ�$�Sʗ��?�wo���٧�6�:���\A���r�e
XIބ��:籾QE���h���Q'�3��<B;C��E���G���|lW�^���;����R�H���m��7���b��W6ho#��_�ڈVw�16?���/3��F /�2�&��H0 C�E`��j����?U�s���OۿO�����(�Kx����H��y(a������g�~�@W�\ўD�ߩ��aOS�Ӛ�^R/���)�T2ʹ��I6�H�y��`ftI��o�}��� ]Ο�62���KO]d�J`_�`��2�����g���_g 4)����}ĆFU��>�O$�?��{�����n?��N
����P}����x�=�fq�2�A�$��=���BqZ��I]� ���d�G��WN�p$�&��QKW��С�N��T�(SN����qz4Pq�f&��)	�q�?�?���R�E�B������賟F��ӡX!�u��v�y�8M.���½� AiN�݈��K��.A�j����Ɏz��/LpV��V3���(,����(��:<�6<6����X�[�:c��'е ?�/�"���h;E��1�ײ����4���\��]4R�ss�\�h��	��cp��[q�5�^Ob�
s�.<S��ZM�1�4�҉Sڃ����k�trREzq���uK�/��N��/�GRvR�i�AI���S��ҫ"+NXzo�!� �Ȩ�ܹ��|-@��-+`��+X������9�f�<!��	y�O�ܖ����.Ӡ߫YV����5�)�=�`��1�+9�OQ����G>7 j=�kg���>������9�&�Ʒ~��UĆ	���'����:��n���XF�� (�}.Ǆ��c�ȵ�wj�侳p�EGt/y�N�&�Ղ��:�����7`7YP��U0�auiϬ�g�R-�`��d�YLL.���A��J0����������!��+i���U�e���ο%�He�V�P*}����	 �~K�&m-J�" Az0k*+6�h6:�~+�}�l���|N��|!��x��5��s%#�|HR- Q90	2�~G�^�!QB�=!�-ã��,��i�j&�=��������Jʻ&D۲������.�`�"��ǅU����&��uo6K�dMO�j�֭;x�'��}a�Qxh�UR�B,`�G�h�y�g_���η���?�����7���Y�^���O#���ի/PZyu~����e��Hn���3��P+JI���8@���P̎O|�x��7T}bj~�g��@`J�\��D�F���s� ��D�_�N�RK�I��=Caj�w��^5虽L�s}�r����GP��c�O|��ħ��|�����G?�y���"}���N[���P˗��vL����)m���̎q<q�s��r�e<r���<��V�舊
��Z���|>���O<�{k)�M��3�����{˪S|��C�X�\A��H��׾lqH-�z�}�����1��;��F��vC3x��ݢYt`tb�<������3�϶;����KU����<�|h���v����J�8�@����[�]��)���h����O�Qbp��j�g����?�W�D>��|f��*}aE�����Bx��#1m�j�*E&U+XTg&��$>�s��{�?�YF2�#>x|����x���F���5�f�����4������YG�,�d-Sr.'��I�����z�L�=6�<@.ͺI/�E�����8�d��1X�0�Lm'0�\�QE��e��S�d�6���1B���4Xڿ����ag��f�
�D�@��y��YJ��k�
YĂn�#�а��U1��+�1�ms���ZoGiiL�=ymJ&�����P�k���1��P{jjZ��̉t)l]C����j)�`�w�ֵ�hbk�J�9�����!A���	��d��8��6�y�*��4�M������`�9�>�Ur�nvjI��5��d�LCWp�����8Pΐ�[�mjօ�0�ξX[	s�PBH��dhL�����#�뫌��'�4�#����d�F�n%��+��Ƈrp����?"���}�.�{@BJ~[��!�M�y�&�	�fyy�W�q��>�"N�9���RJ�������T�{ ����I�E�O�mlc<�S�K_l���+0ɞ(�Q)���0�>�z���\�G�lC���R�D@�n�Lӳs�}�
&�F�~�X�uW%�:m:��� 5�5h���^n�K��]ڠ��\1P2r�D�%p�4P���p;�����[�]�XO��j��̓��]�a~i�t	�����W�@���ViB���s��I�5�l��؄�8௿��W���L GBQ���
qrr_�!�^�Kg._D���K���1m2����{������������A�]:�f��,R�^�o@�ͽ%*2�.����f�.\xD˽��
xz�gp��--�sD;Y��^^K>���絜- �ܹsh0`��D��褸�ܿ�@���ٳ�!ZXX�}�����r=�x�/-������{�ï����փ�P:���~���� ?�^c��2������|��� >��G`s���o|���HN�I�:v�������G:���5��ӌtي�N�\Iᓟ��~�3�R��/���X��!WJ���ʝk�Zx�F��Ao|�>�)��ʏp��I�6�N���!8�m�����_�%XB�(5=����`1��㗆P�����wT���HX��3�c�R�F�
s����?��)����*�g�\�������Xm���B�����2��~�~�gdL��l<w�b��hQ0�3t<<�nQ]�q��[j��Z��혝9���bS�^ć<<rU1�LJy]&�����X��#Q7���o�������Y�2���x����*��\���6�Qk�p���ݼyQ�&�o��@�93�U��_�7Hn<@�~���b��r���w����q�A�a�J�Εj������,s�oB<>x�����[���;:-)ri��ƺ:)5	0��ȸd	M�A�ڸ[��i�GL�42�4��-�y���R�H�'ѐ�F�D� b��(�?F���5��^b���ƶJ��L��~�P�/�N.3���?�#,̍b?��:A�3O<���}�Q,�}/��U�63ꥬ��=� �tģ5"���.䋈LOt��+W��eU)�遼��]�鐋�v�U��a��ᓞ-�P�عt�x�x���c�]��/��r�f�����3/"C����kp�-8�-�8c/�I��4#��/�&��)�4�� ���������;o��5,L�F1[R9:���2Z^鶤w��e^�=�Y�ڇ$�Lp,����:h�J%�\Z���ӆ���C�;}�'vn����:=,z��$�4�"Qh��"�~��P׫��G����Ķf���T*�C2E~I{��w�x��m���6�飏,*	���!�G��U��O3Pi�5ܪ:����$���6ׯ�����Ic��B�%�m-�_Y��_z<�L��?����au~�:�ܗ�We4;Ul���'��cS���x��YiÃ�����Y��5��9�ܯ6~��AQ��lt$�{���9v�v-9��+�Ut;f��.g�כA)+��w^�1�cO j�|4p��X�V�������t*O�8��u:��R���/)�
��.e�b>;,!�	(l��k��j(bH�DΡ�E)�!?��\hil������*�pÈ�����K&DK�<�һ'�2Q{ g�4�,Br2���{!�t����<y��)IO�L���������T�/P��ͦ���deOI�!�����^�^�+��i9O�٣��ejY�e뀔�)�
��@ȋ�4���^{�UL�����`{��F�}t��?�R�g���d�Ul%v���&g�xn\x�n�������1�Ơ*#�>h��]̀ʚt��:u�'��������eL3��۫[|.����0�w�y�rZ'P7E�6}�Y(2�@sa׼�Cj�{�w��r~��mt+���a��h#8,�.Ҽolm�s?[�Zm��#�UZ(3�t۽ʍW��a$��6v����\�Z#��4�a����)}#����P<��z��Գ</=ma���B f����5�����IxmԷ�w:?�K��v cؕ:n�I�����G�A����32\������ܧN&����d���GH6��㵗{x��sܻ��1��~��hH�A����'MU�C8yr���_���kڞ$���."6�n�A�-<��.}�	���
x�3`g���>�Uzu~a
��ד6�SS�j��`s�N����6��>�(�5�&��##1;�BA�0�p54(aksE�4�K�Q��(w(Ef�C�==�4
�o�gd:E'6�]F���<d"�E#e��jA��� �-V� J��Ap%��"�me�*Ӭ�4�"�C|��"���B`ؠ����q��+��'>���uc�K�㑋� K�����A"�E���RsG�M*K4�Ui#ɞ��Z��.D>���Kd�#����^�7Asx�4ʍ&������?@>��I���ьf�,��t�F*H#c��=�sA�s:�:j��h�@����W���!�ar ��`�k�}02�<����)(Y/�m WVo�035�{����s�!�Ã�|�X��m5	���YV�<�X���ڀTZ&c�&%Lղ.A�!��4|�k:2?����b<���N�I��?���S"#�%k(��b��jx�\����3x�ɧ෻T�Abvv6�������_�5Ć�q��YLܫ����c�m�l�Y|33�x���8�D5�*�A�mҁ�{i����b>G�N�����{= �NO$��%R���H��!��	�Wh_�x�ի��$�w>��i$�`��T��F��>!k���#b?/���}#+���wm�{2�i���3�s�GQ�t�ͽ��?E�[o ����J��������Ȱ�C�~C�:� #�W�0$�'��IFP���n%�+{�\���D��Pņ�
���K9N�)J�%$�����XӒ��HFO2��ݔ�
�Q�Qh(��aS˵B�$�i�^��p�
7��A���d��fuT���/"A nbe	\��zS�A��n45����P95�6���E
���	�m���Fjd�Y(�F~2u/*-B}"��`���_�u����������k��HԎH|ګ��U^7�c����	��ӆ8e���:���X����)�ʗ��v��o}�A�8�����S�~�~���_��W�3M͍k���(y��Ɇ�cg	:��"h�д�݇������k��+��9�����/�	�#�����`��&�|嵯cm7��|�o��'>�ja�ͫ�ʿ��������uU��F s��k��� ����,��w�=���Q��
x�?�Af'�:����B�C�]���M�,0@�2��]{��/�C�'����U^�~��v�V� ���_p$����v���ǁr�������i>������`u�0�$2;�`��`��,�pH{�Z�������;�P�Oc��c�{��oa�{)�?��4���Y���X~�_�����f�e߾u�=�Ɔ}��k�ٟ�	B~'���$�x�eX\�ڢf��>�x���ٳ繎\�7;��G{\R5+Ѯ[�u���������}>�w�X&BU�K{�<��&�����ظ6��h�<���8����y��>,.N!��ad�B��Ľ�GK��mFH^;�'����!+)!�D�2�h4�l��F����b��ƹת* �#���cH��@�*e��~�{�������y������;�y��"��t�I���[Wn#�����yF�9-���|�;��[��7vpv��W�dضw2�~s~�/��'���������f�ş^ct��IX�����0Kۨ|R^��ZV��˛p�nc��.�C�a����?������������mu�����M�G�%$�.���W�ّ�.�S~��ݭ������٠�í�QɃ%k'�Y����ԝ�R��v�E[d�@�,��b��l�qHߛD�q� )OJ)Y�V:}�.@��{'�!M���(A���9ү���J��L�on�+x��o��L �4X5�x��W��f���+��A��!�㓳��/�Iy!���h'rh�Ч�,����,*S���ӓ8=���^�N���(�lN��ۏL9�
j>kC0�5g�&D�W��8��gO��w^!�\��g��02E���e3�� |t"::��?��an:V�͏C��|�{.bӾ�A��NM��v���lڔl�j�ƫ�|c� ���4um|��մ�+yȺoo%�^gAћ�r�����	��`�=�s��i�>ɺ� �dw�8��O2� 
���KQ�0�$fC��-Q�=)�/�_2rG��"+'"�<���uөK�����������?�q��+�W��:]}�#}Z����5�w0����-��'G�������7�HT��\���|&!P��������1LN��5U-<E������6��],Ny��-"���'�/��[�F�\�|?���� Z�R&�3'��b���~�jׄ�3��~��k:��s��Eڲ{�� ҡg�(m<4�f�WI�S�*�]M�M����[�����?�O��S�Ľwn❻�<����]�Ј��Ʀ���}���!��,ϝ���{7O3@;O��[o\S�ګ�Q�M6 ��M/,�38	�l �����-�~��pyK8����x���=8�v؂È�Gp�UG�dbй���}�I��A�~d	w/o�~H����7�q@�/=�2̥,
}����+���q���p���jO{��ս�o�s��J�������8�Fd���o���2�G+���oea�ݖ�J�MEi��m^�&��'�����Vj�"��K8}�4�t�o]�ڊ"O���D��d�K�2�?v�F׮��]<���q�������VD����5��U�3�(���￧�`�S�����7�]nV'Z��B;��#{ؠQ�X����J�Q����2�ԙ����(��Zo�҅����4N�4�s��e��� ��tb2x��J�P�SDY���4
g�����ӳ��'�1O�K?�E�L�����e����:�[ x]�?E`YG&}���_F(��_����Fi��^�8w�~B�ۣ�����34�����E�5�x8���4Bޘ�#��U|�S�F�8���g���f7�쭴����t��&�g�S'}fwo�F�^��]��ņ��^EzW�MN;cĊ���km$�K��\���'=�w��q��i܊��Q���W�.�@8^�w:=:J�ٔ�F�,D�>��|H?�8���z��l�/+�o%:��(��|`�8P� ��L��8�8vLA���
8.K�q��"�^J7�9U�L�	��K���i����/c�A���qv�@�{�;��*��4p߸��C���1���;J.-�����Gx��<r%��:6	D��wv��S��F���T��*�AT|��<�/�#ͽ!0�m�ƹV�CFE��Uc��<���e宫��r��o��_ ����n��F$lC��v��=:�f����C�?���=G�QB2��Ȑ.:�T��Lр��2j]#޽�B�n�v�{�#X������Bb���-9O2X"�~��	��{��Z��d�2n>%�j��Q�LM��&�}�x\��� A���ʰ� Ai=0�*m(|��\�C����V)�;v⽒���GU�30z�����2	x�<]��d@�Ȭ�$-���)gK��d7%� x�ʅ����Ԏ�Op�D�gY*Bo��H��z�ʊ��
œ��r��@���r�����p��eLL��D�i�+�	��ׅ�D��A�.cご��RE�j��~׮�E,<��.���w�NV����]���{!�Y*V�fJ+`�-,���s���1��:�n�x����Ю��������a�S@���a���T3M���{R�'QM%p��}̍�����8Q���E�x�;��̀�������;�.���!mq��Ș�5X"�0����=�`(�����Qlmc�Ab�A���c��x���i+�]I*Ǧ���}�t�XS3�\+�[R���F�� _��_R4���Y�_��k����[Q[�����U�.�d��#����N��x��<��r�'�vwQ�I��}�ǰ��� ��?6O�c�*_gjx��v��a�w��5�c���,_�����U��0<���14�#����Mܺs��o�<>񱟁��}��=�<�������=�`)O�N�`�o������lIO�UE�f��;�(��<<�mf0Yz�a�Ҩct�l�	IZ&0��g��뛯�AOo__Ǳ�0��BL�D�®)~�dP�&��h�xZ��=~�O�a>�b/[���Hߋ���_\�4�Ns~�Ѷ//��1��3�t"�HT&|�'��t�.ܧ�6�\� 0ť�۸����-«E���?��Ȩ�/W�9�s%�Ku�!�
~��@0��k�A�Ց�����@i��(C�6�n�_K����=�[��9���m����թ�R׀W[�x��GY%`�ʿ���L����s���l2���-���57L'�rZr	Z�/G&��{<5��؀GP$��1�f�%�U`^,
��>��+y����M /�VJ��'N"�!��dS���/_��G/(7��Ǝn+q�GZ�ʸ��.�C�5ч�+A�ݛw��z0��!T
)�*iܻs����k��lU4�iW� ���{w�R�����ʃM�*7�Xݸ1 �v� @xf~���a�:(��(��ɓ��}��:�Y���/p��5�X�%��ذw�*_�A�!r�/������>N=�i�������?���:v6�j,�i� �0az��:�b��3_ȍ�o"��aaz���_��B�a��gat���0�`l;i��yWn<@Oh�xv���T>:U'�d�󞮱d*8�t-l����l--1�D�I��r
(let2���8qB�L+W�k�J|��P'��t8*�tԙM��^�$Ӯ%�N���S`�n��
Д
�`0ɢ�Q���� V�0��B���J�?WWW�:08�~�u���y_Y��GW[&l���y=�K���*�#
�i"��1:4�Xȋ`ċ���6R��C�y>[]��zK�R;|�#��HQ�"g�k�f09>�+׮��gF�����7~�o#h6��w����ۗi7lڂ��M�̅���B&W`�R^�jIXU��lna}�F�~�����g/=�$���y���g�?Ԁ��6F<��]�����W����]��m�g?��Ņ���u�,����H"u�� ̍tzOě+�h׍�\4}�"E�d��q���.:;i�.���{w01���7na��#0�-e���yqw7����a���yO�#
����"P�RQK����G
4q�;m���y,z�Z(#��#`,�� %�x���_�*�0U������ʯ+�M	6V���
����R�X\�w[K�6�3/U3��@F|���Wq��������Q3�G���J��(���i�K�">��0����ku,;�����B��9H�c�2P5�d��l������|�/P8��6M�*�H��3��g��S~9��)0[�Uc�Z�bm�ȃ�����+���+:m8?S�sO���s���+�MݡQ��̘#!m�Q��:�*]H�*[(�Z�J�IO[M�����'2-\m:�����������?�b��n��`'���!XZ:�$�A/�4:&9h��$��J�hG��H�i��>D�$ϓ��
:-��6h)Y\�,��K�����~�:���@���Xgzf"%�n��Sv-:�ی�3���tl�4b�W;�!������4�v���M��vsP�m�@�e�0���٠�)���IC~N������u���K)���j�L�4��>D-�q=�(\�����b8S��uX����M�'���s��U��K�����1�C������!z�f�;��2AG��G���I�r��$&;����������?oc�`eLR��6��HW���xWa0�4c"YI;],Ձ�\��p1I qr���\a �ϵ4���\��]k�ʸhrl��̢ӊ��1��������֍����x��g�ZŃmm#�������=�MΈ�vw6�#���m(>��T|��.�u=*yhro��3(h�ajc=��z:��%:�<��Q�ΝF�oǬ׏D����{��I�~�6:|[�?'Q��p
 ������ө}a��5��|:�ed?Б��du؄�[��nܸ�=��?(C5R�������,�A�����5(�t~��|Dt-��C��_�\��o��"|i�w�Q����T�m	^$�'�VhcP%�{J�-Ғr����U��s���uߊܠ�=U����̶�k�)�=���:�����bԇ���/2 �3�����x=1�C�*�lo'�|C�4y/^���|�:?��!��[��g�~�����;���7���P
-,�����B�N�>����x؊D���k/�,U�4��ag�Ɔ�񭗾�K/����"GP��D_�L\8x��-��	8�Npp��l݁+Π����an�6ʌ�Ǘ��E�\��h4�wo2�	�ab ^�o�G�4<1W8�ۛ{h�M�,����.z������vx�\� \�س��y���P���JIJ�*��XL��-m;�R���A�P�B����cvj/�r���d�6�I{���������U�.�Z����Y(V��1��-�O��4�(��b�g����%��R}_mi�v��h�E)%�v��\64+9���Q��ZL�T߸�_�ZD�������p�
l�⣣�v�ZI�h��޲[�HY�������)�����z�Ka�Fel�:i�Q����6������{wua����x��2�>��s��_�M|���s$߅=[�����01¤#�����8�ci8��>%1n��t&Y����h���X��:��.U�a1\�W��O14s��Ӥ!��H�a������uf2yH��+HB�4ߋVo^�$�z��f��:�D�"�+_:D�N����c;��F-��~���;����a :��]��,�Yԅ�Ɵ32o��\&��*��F��xlj+k"ᶎS�N�ܾuӳ4��*�%����	�t*e4��X�(�k��)f3�Ԏ�CR*'(N^�qr�W+�;&=XbxEAB��Z]X�Ҿ-�6U��bw/�����8<v�v)ᔕ�ߩ�/W(*��d^ښQ�����L��ȼ�k��`P�������&�T'[���;��2�>;����V��#�8E~���c��!Db(�vy/y���{yT�*M!P�+�0�}?��G�sk�.��˯���S�8��c(�!���<=���T0����E�o���7�T��c�����	��s�\�$F�/�E��o����.�J|ݪ
�;�,���/��j�W�"�}�C��{�i��v�U�s�^��$��cdw�:�'y�	L-^���	L/^��o-�_�6_߂8�G�*�N�!���F�[�=!�O�jˑ�F��2�+T-�19j58T�i8(��(��}!ϑ�
0T�g���k����$k�5s(�U�-t1��l�>��I���4� I�Vs���z���}UyG$��c�A�/�n����T�wB�3(W������wr-�>�Yd�DyF2�3J�h5�����z���Sg��Ѭ�s�J�_�CL����4�)�Aj���?�ǿ����1��k@-�()���-�M�����^�~�F��p���~��m���S�;!�_[}�=4�Ӱ�'�L�u����*��Bxr���+,��׿��g>�]�p�J;�h�Wv��^��	�������ϕ��h���, �ęSB�m��B u��ծݓKg��Y��3X�}������ǰ��mr��=F��Nb��UL��҆��?�i��,.�B4������,���A�U�=��6�c��f;1�(�xo�p3�m�m��N���u@�ޭkx�����a���Z�d-��T��P���3���x�9[%���Q/�m���b�/r�U�v�Ղ��E�^�2r���_�-w�'������h1��I��@�.}��9m���	b/�����}ڨppY�f��ɉ!�C�����Q�:�S�xߏ�
S��AX_��G�}���hm~�8/7,��	cnLΜ��ڂ�݃�!"vbjv
.����1r+��S�[oQ�la=��d$���q�5�M8}x E��Pn)@4`��SG�F�H��;��K��h"js��ٳ������؆�*B��MF���mt^{Z���n!cv�vi�E��C�������b�tde:2F��c��Z���р��E�f��K������?�3GL�8HmiO��#T.bp�!�g]�%^X"}�gDz���a:�1,��a%(�!W�a�я"�����}|�;����(�ڪ{��
���:���\�k��8�ݝ���C��f��/EJ��1_����L&�s�2�)�����9��Z���tJ�AiYA�d(����H��۬��Sڃh���Õi[���pme�4(��}0)-eA�ӭ�J�w�Y+�7R�����L��m�$��E(�5�F^�C�)�'�E<>���=��lwJ\g3���x'����R�ar� {gO��;*���������vS����f+�]��#�V�*<L�U���VI��n����1>��+ ��~�p��g�&��W{0��(61���=F'<Jg�M��ɳ���60b���)�G?�>���"�#�(5�x��&f�����������C�G�H$w�Hmc��3x��eޣ ��!�K���b�,� yɨ��0|-�Jy~NN;
օ�Y��L�Ki�������(�H�����J"8�% Oe�(����R�%�O�Cʲ��xt c(�g�A�eHE89%711���AY�+Y�a4i2����󓲮P �>���r$�O�� ]��ՀD��epE���|/dד��x��7q��E�;;�|ݬf�����r��x��F#�P&Io0?C�d�a"�Ǌ�[�����/��,���e�`mM:�~���!J�*��V�)��giff��_����%$vӸv�&��%������!�z��VT�cx*
J��<R�m�۴K���-��]�,����Gq��)��(1��� ��9����gm�;iE6]�n���U���E5WC|x
[k	�?y��S�b��V#���Q�|_"��%Ѣ�9�'��i�q��*N,�)�̮1��������;7Li����<���l|�~^�B�����m�ݫ-����?6�l �j$2l� �D�(�]���Ȱ�D��^$,ОZ膤�T���v��w�4�>P^>�f��~��O�"$�BX�6ҫ�4;.լ:��׎Z=�܆|�pЇN%Š����q�7_E,���(_d�v��#�k��02��5�8yNK��.��|�s�gf�搯;pw����1��m^>HZ�����|��A����+f�/z6:�.jU#��uB7{�g����vN�G����M�({~����B�5�r��;��q��,���_��S�<��*Fm�;=(R
�|�6�e:���{�<
NX{F�Ǎ��7��Mƣ�*"6T����m�rq�����b֔� ���k
�\76v�ԡH���S4.t��&��� K{��o��cQ:�;`w�NnV{��g��l5���ѢH����h����~�n/���#[2hpe���gt���s��=��,�ޙc�`|b�q\�qEK��
�/���qh�����C�,��d2�3�	����Q������
x<Z�IF� ��C�)Yq�Rv�8s��\[�NK_��n����3(9KfP@�dl��Nx�j$K�NH%C$z��OU;d8n��(��L�J��72�)�SJ�6����b�*-������h��J� �Õ�p���i�������?�g���\�p�I:aCO�{��ǈ���p'�Hq�[f���` �F���=��X��R ��>Ε�P�s�ӡ-��;8��E:�QD'���_�:SԎLv.�5���O����1:^����(���co�6�{��|pI[�ʖ������1t����k9��:h��u���w鐄�0�4�TdЫ�4`f~�kSQ�N!lvD�z��ft���6��TְN0���B-��G����ޑ2Ϳ�hj�_�{I��d��%�=V!0�)z�	��3gμ����3??O����3��S:#<���,�#|�`e�J0#$�G��Bt~4|rą)�E铔U)?�>���uKIpl|�֭����->�ߣ�C��m����xPi�dMR�=ܼ}�A` 1����������xu:���$蝡h�֝�p�	�ӎ�X��2t� ���H��&�������X��s����M��F��_��"�-J!U�z�ܹǵ�"@p�c@�	Ok��XC�hg��=9��;�hw���	�Ƈ	�Rp�]�LmUvʕ������J~�������U� ĳ�&8�J��mD���;W���	(�����Y�f�|6+����d���� �"�A�}�2�F���6�>�o,��3�p��U��7F�b|�������V_�Gm1h�7is۪�c�B}���&@���䅙gX$V��&��;�Q#��䶹0��%����!�H�Vpl.�=�&3�^����ǧ�V�i\�������r���hK���Y���V�C_$k���D���#Y�"��q�&��v�c�a%��Љ���g�\�u�+�WU/g�!g���Nj��@��%�#�^�f4k<��x�l�����֌���l٦�mi��(��l�)�nv�42���c���}�=�����j=�zU�޺����'�#=�Η��DW4NG�zt=�Z/eN�[V�1�}�q���O���O
����[zBJ��b�%P"̩��0�0��Q�|�^g>z=���B�N���h�ޝ��yS�m,p������|/|��^���M���7�@E�|� 6��4�e��!*ރȧ�h`{�akҠ���~�`c~/��GU����T*C�Dx��7o����׾���.����aj�2AZ��c����,�0�ZhQɋ�c4la�L�>n�Xįߺ���?�+o�����[=ܻ�����sA��MĨ�:=��Ỏ{�G�A#�ޥ��G��! ]@���������wq��G����4�8r�ƍ�����m�ޗ~'�Ƨ?�ӆ�/���4�]�Ǎ������[�l��j5�P���}�U����;��PC�PZ�T�Y��@ZQ�}�(ba����;E�M(���EU'���fsk8Z*f����� �x"y�t	uF+��o��1�C��"�R� ���|�s�é�'Ѫ�\4
����
��Q|����g�����ⲥ�n߾���^1�0:6C�_G~�2.��t>����I�bym7�a��M��mU�7:6I��u	��2���@�%�q�Q���H��M ���A|� R�)�m�J�Yv�ҭZ:�Y�aqe��]�K݈��a�`l{s�ܴ�-l.�a��~tv�΄�S�h��HB�0z�=n�B��)����8r�e�]��^)Y�0M�Mc��?b�Zj �Z��Xi���`ee	
#��O��[�nY3��x;�M���x�tZ�,�l�'�D�VV��I��v*E���G(��L�j����+B���e�Fݽ��0��E�FGFy/7��O`�s���`2�5����>�9��
d�5E5_{���79z]��"Җ�K�Uk�Ni�*uH�;�����I��&y���E�_�Ћ��7�����6�]��zyaM�YY��ĸ�i�Gf��{8z��޹N�Q�3��Q��a\iy�a����`�%j�(�V������a���{o�g�g�fG(�I:49\}�2����&��q��:�Q���}7�\�t��DE�U���H�	V���Y�L^�S�Q�C��MCi7*H�Q�7r����鼴�ۖC�>�Aͧ�A������E��C!s�ݸ�!_.���R��7����g1N4���5\S�ki��6b��;y�Ԋ�{t��^�I����U4vј��X��m�j���sS��mQ��9F�����JX��tafg�j��ɶ�����?�\��uR��t�C^Ĺ�k+8{�(�/R�2�n��,uA�İM��a<�W�SF�ߴ�P��1NZ]�Ps3C\��e���s<\�E6W�
��q:�1���Vo@�O}��wmoz�=��|�&�j�iM��㉏'�N�WͿnQ�Dc!3�ݮ�F��!�F��tR�+�$\|��6�(f��T����;���(�����y�Ӫ$Zn��C������U���Q�_�sqz�3���@'�!,m��c����Ae�*����W�'�K� &�B5�cms�<��&F�Ʊ��B�Z��P���6TS���wr(��.�����yden���"��5i4��a��4�����=̌E�.'�v���ɍǓ��2%�;�<&'g������}c����.!�	ѻ��ʵ��p��W��,�b
��"@��봭۷��HgΣQ� �*e�RXJը����a|�;߳�%}*��
�������Ҫ��~��-��x�G����){�R.e2�2�*~���`f�ޫC�E�T/9<�0Чi2�Z+�U���6�Yרךf�8e���b��͖u���׹4\t��,������x�rQ�~y�����g>�S8s���f�а�q��E�#���C`��A��a�,���kX��FgP?7DcTl6���Ӷ^��E��r��[�?|�NA����P{��.�a��8o�{���$.������Cr.��Hr�|��!����5��j-O���� ��Fpf~_����	>�����6�����Zt5Y�e��S'���J҉"�(}ք?A�R�/�3gN�;�䭶��y��uQ�����q���V�-<�{VS��"(����,Ф�|[��)Z�H�Ҽ:��>=3e\n�]�0F�6�M�`	�J�����ީS�L>4aB�"�#e�w~�w(�qKk��!�4��!��c d�U�j�Ųݧ"��:�G��J�����P[�i=u��H��S$�&_����<�>2nΥ��tt'����wW�C=���~�S?7�hf��-`bl��?�G��"����{o��٦�<��w6���zhҘ	D�� ��$��N$ba:�ԕ&3�q��o!u�?v	�B
�c�tj�(�x��~�]����x(��ϟ!��"�^���<R�`��`sۡ�k����C�3��t���z��87�w2�^���H��s�P(�Ys�3t��1`�����24n�=�&�?���4���fǱ���u�a��V��[t_ZH7�|lA4�N����4֗ބ�י�.�) ��9�tیCS��g�������%r�ɳ�_Rkz�&9��X��u�k"������5�Z9اN����u���(޺z�:����V��2tL� ��Mi����'*5����Q������"�����|��ǧ��!�L��iS���d��'���-~�V�����O���xz<��Ġ����m�����
, _o�@/wb� V���!Dc�
wQm��Oݥי�椡Fv���1��y�\E�E��tN=�������[8z�4F��Vw�i��4�IL&h�����j�E��M��^G�7��s�⍫��dƩ!�8l��]x�.�d���G��C�G�,8lFI�Y�ܘ׷U� ���-��ͻ�ȋ197��~�ppve�CQ1�.Q���vX��#/�o���@$6
W)�J&�*��(7x��M�Ѯ]��X��}m�=>�J�,���ȪR�hlz�N��nGO_�������5%�B�r�54��%�JZ�������"D"��|V�52��u��-���7+�h͏u{"��zl���RjO���$�F��ֹ̦�A)�i`��ppR���UP�T��1�O���5�\"�1P�&���i(����6��G����@�	D�)�]*�����~���c<s�E���?���x�T�����W�W~�@p��e�����Q��縊���4�;�~ui���F\�ull��O�O��9�w��Z.�-�P>�꼎���	�UW6r���N.�C��v]�����v��#]�)����):0�k˘�E� �Z5�N^+E[�96��P�����4fch9�hx&����`���޸��thj���[���3�C0�p�=sM�mmt|�R�Z��p���\ J��v�1�S�E�N�� ��:�sV_)��N^Ec�U>��9[��P�@��v�;5�$�����m��2^9�ӣ�E��# (�����,/�82<�{(�R��D�N�A�#R�X߲�)�٭����9�1��(�Z�hE��9�LvPg�$PÓ�95=a�!��wP[�����*��Z�F4�ËϜE��3%e�՟�1��?��k88����8W�Ƴ/�(�G��������/W�|��m|}�
�Eߦ@��B~{^�g��v G`�C9����T��/]|.��kz�d��C���w��n����������qkH�fwpxz�Z��]�JM�63D�'��������UA��~��8��pj.�w������N��יN��kc�l�b��K������s��ܻ}�:�g����Qu������±��`$�E���Pw��s���3&�Jw��"����7E�.�Z�2����hW�ǭƞ�ꫬ��1��,��J���|����@Տ��(�~��4��I�WW<�!�>jռ��(�ڧc���q/.-os�m۞�z�$�E[Jyd�:�^F2�f �IW����v�6��Sں��ӏ;/��tr<G��~Yhs�e���e�{]��ɼ�w��6��~O]}O���O
�8���qgpC�D@�|��q��UEO#�G��O���C����4Kw1���}E�!lo<�g4L�Є�T��j�,:���H�����ݝE��L[]W�o�:U��2
Q�ȠY7c[`5���B2L�І��h|d��2B}n�]Grv�����
ȓ1D�#p���I�,�"�&�Z~���'�azl���k��W�+7�?Gbx�|��n�F��#6��@j�KO�/V��q�u���/,M��ͷ��&��³'���č[�p��q<��Ʒ��GF'ТB~����z�<|��T�z4�S���VvW�6��;���%�.��w��i������6!���0kvf��2NP����	ZJ����x�J�j��#�葀[�V4 )c�)%z�:����_;21f�u����* ������E
=�%��� h�������xU%��Sg�(����������x�+�C�P����C\}�-L4�)�Ư�3�/D��1
�^{��=��������p���&�9D �1����EYZ��)�"q>'ѯ�6�V>1�P' ���7�୫�&����n�w�i;j"��7*F���,�:�0��� hBÕ+71��r�~l؞�8;e�h3A�C�A���B�L�B�[�zh\��\}��O�t����?��u�6��Uъ���:�T��E��e�mM�ZP'f���^�f����x,�L^���x\^^2�����l�4`D謴���w84�VN��/��C��s�魨��Ӻ��u�m��v�rBt~M�Q�����U��T$��¬����n�c9u��O�6!6V�1kʈfs�z-�/E�U� :�Tz�8�b�O9;���N��~��[J�Qߤ�4�����<7��f��L��¼p�<.<���Vp��;��th;��	곶&�L#:4���� �<M=SB���&�Dd�ts��|�5��.D)��a��A��1<{�E��z"~�$xbAl���s5	���l�"�l 0��N|�r]j��$7��-�H��bM��-:p�y�戾�s����-�#�������g�x-}~�[��C��Qu�f����D�J����l����(��D(�(7��SnL�ƕ&b�E�BA'�_�:q���C�ac]pRv�!��:x-�Q�i�ۧ���6(F`�}!��^��C�n�2;�]�R��%��w[�q�^��Y�-�#�/��N&O�$���9�]�0E�:�0�-�5���n�7�$#٦]Pǹ	�Zm�;m,��@��N9g3ﳭ"Pޟ_�T�=��h�&�Vʔ)�����§�OXS�5ħ�)q���Z�p j���V�O��b.�/
���K]�.m�@�Jv�e�<% �F+OV�&����rWqn��B�Pk)T?A��<D`�q$Р����hӨyЃ�jDF�]DG�ȍ<�г~�+-8{I�yw`}��S'>���P	t�c��i<x��_��?G� ��~���衣����*~�K`�>��Wi\F�'_�/���ǟ�kt/��?�KT�<?�'O\޻�^��p�"v�6��m���j��|��:Y	���YW�?Aq=��^��m�ui�5c�[>F�Zx��;��@+wע.-:���$�hQم�ݹFa~(D������m҄�v��s��O�5��W18��:��ۣ�1Kåw	���0j��F����tP��2e*�,�_��]�i��v�@��f��H+��$�a���%GFr��A�S�w��p�ND�rT�+�,�k����ｉ��+��3��Q��Y�}�$���$nݼa�qv,�v�>.>;G�q�����t$�U1W1�*�(q��GS�]�ǵZ��#��bz���O"|��[)�f�Vq���o��-�=�h+��N�k+U�1�k�t������j���3���e�Jp���n��M$B��y�!x:M���Og�.4h�H�H,1��
��8����bscގ׺�=�څ^^r(f�F��!^��L�iu��x�f�F��K�΂\���O<��'�e��X�������q`�T&�W�w:�j��l��Ym�~=�j�$#�N���.��<�ܳ�>��w�k3�E+$���7_�g?�Y�M��ڵk�Ј_���t�������Ţ�ϗ���������h�G9Z�͍5L����G�"1�����#|�?���Y>� ��z��5��g~��U�ic��A���A:hD>\��c82M��#����ء�I���ab� vv�V�;Aݣzb��ON��sD�'��N9<s�/q�w�<Be�m�6.�H���t��;Ȧ���v� �N�:	L�Z�,��\�RlpU	>	��5�	�K��:��h�EGIM�F���8m�de�j�=y�6�<x�r�z�z�μ�e�C}������-�Ю�Р���a���~����h�|�Z���I.d�����(jM��j��^���������צO8��={��ཷmrV[�K�Y
v�������h�ɪW3��h�vv�n6�0��$��l����D�n���?��M�t�NJkա>�SW:42��ҥ���;:k��]����ɺ�Ak�j5�;�M��Nǲ�Hr��;��E��Ձ����	�'��~��p�,D���&m�k>G9k]��>�"j2�
gN�Żo���{q��Bn��=��|]�)$�cƳ�Q�� 7P�^g�J�Ie��;���`4�D0��$�C�֣�N˰u�*J��:�����;�x������.������_B�w�v��i?�#?i��"�9	J�~��?��.^���O��$��/��/�̙3x���o����ϼ��11E�K�����_�E������$?�{h�����U���n����o���Ib+L���q2f�e�zxu*��ك�=�6U4�Dl�ưnJ!��ɠ�G,���Ћ% IS�z�;6���,��gf�����4Rγ3����!CX�uQo�������k/uo���5`�g<5u��H��S�j���C܋�F�A��R�
j����w�e5�2λ�n�ʘ��>�YEE�]�~^__\����qUj���f�v�7�*�^J�-A���V�hC:-��Q��0���h����:�ﳍj��X"�]>��vN���K��A�K�]& t��h��\���L��86l��S�����W����;ІiV��ᅣ�0����i>����W&��	�fn����7c���*V6��E�+���Ȗ�4^"�w��%����=��Q���k_�ц��v(�	�U���s�Et�F��&#�u���g.�]=k���ɨ%�y��ߵ��	ti�i�S`$ϔ�R������J�[�H�Ί �A���P�O _粆$ʜί� ����t^�G�0==m+�	h
�^�~��t/�`���v�����h��S2��p��{v?�Q��_�u|�cÃ�-�����1K�����a�P�����5�Ǉ�(������ud�0�7׭�X{��Y�\�y\8~����{_���sXy�:�S>���wxf�kK8<;�O��+���.�e�d�r��D�Y��|5[����8� ��f�z$��<Av�X��Cg�^�<5P���`�a:֙,�<^��N������i�f_��]ΐhƄ%��>��G!�z1�Ռ&gIM9�AS�����@Ӻ��p�x�#td"a'���?�_�+��W�$��՛�]���������"g�P���$Az����"�^c	��9/�&�j�m4O�ܮe�j�&���n��ڨ̶MgQ�J�h@kuz�.e���f�o�>M@�|J6�I��?Qu�	��.*�%e���7-���$�Ig��Q���}V9l�SQl�l�{g@�%��3��i�+�ᤎ�5������}4kӹ~o?mF�S3y�E��������� ��Kߦ@��Cu�桡vy=htD9�����ӯ~�#G1|0�;�.cnJ#�T/�ѫ#P(ҳS�u��a�����-������z����Vۊ�E���X��U޻(	d�i5��Pr���s(nfix�4����;��?�!\��6�Q�^��ӣV��A�t�^z_������������o�w�D��B��NMU*�~߇(=5�I|�ۢ�9�ˋ�.�0F&����r�	M���}��8��7k�L���R� /�k?��k>��n;�A�m�a�rtw�!�����(
e�KnY'��{7���O�N/�V�":̵pǰ���J�I B@QB� �Tj{čf����E�T�?t�mlo�����z�P�b|[g�s� ���I��hA1�`:5� #�)���f��P�'�($2_#Cwz�ȴc<� ���%x��""�B�a]�^g��n'U��N	����HN��3"D��6@�1o��~A�[U$�4:�nߺl)�~�k�$g��O�����-�	����*p���T��ʭwR;�8�}0<5��CG�V�c�� ����E`S3Uǥ!@��\Y���.���C�J/�\5M��������p���/|�38��'Q)P߹K��C���݆��n�`́��[�GO���C ���F�m>��83�eP�����}<ED�M�1E��hu|}ܿ��xaa��#�浉0�T��=�a�s(��dT�S�z�wޡ�r��O�?9:�g�k�ݐ�H�9��RH)�&����4�F�#�"u7j��4.Kɴ�%+*��<|䈽_�V��'�/
��~�k&��S�W]�7n�0�Խ�5E�t�V��p?&�������Z� 9��H9^�XXC���9���#���slu�<���G�������'�
Z�U:=���),?�cqh��%4��w/��:�^U�U�t.��s�{qxăN�2�&g�(��q�G�����1ӋK˻�|x�7o`e'��R^Y�Z�{><���Qd�Ct�a:�&9#y��������	NB'6�T�c��u�n��R�xÉ!��؏%�Hm0{;8u����%�U�:�c�xQ����$�����.pv4��g�S�|e:nr�<��BAPj�h��o�x�����.P�iN��*��Z���.�󂞋�9
l)"��@�u������t̥9�n�Ƀ&�F�Ƭ�Z<��}e�$C�H��k���g����1�}Bw��{���￾�4�1P�T �ǛmQ����QS�"��<�>~z<���5�*�!��(V&�ֲ�v�Nm�p��-�N �w�X�{�H����]�����X�0��ݠ�RЦhrԸ�i�;�
;FnKM5�� �Ҍ]񣉈t(>B�g�P����)��S\�"� �cv^<z=�����%�Ζ	�T�V�Cz��,��'-j��Ґ�p|ⓟ�׿�g�ٿ�׍���������W��*�����Uk50"k+z��{�[�M�,��~�V!���A&��n�i����X�JQ�,�����z�����v��(\FYQjћ��@���!�o�k�w�����{��UJr;�A�TE1o�f�jMT+%SZ�eQ��O��@@��u��ј:Er�4�����QZ�V���������oe�Wd�E)��(�ߕ,N8y���2��S�I��R�z��"Ja+r#�Q�Ԍ���k�,�����u���y�һ���dg�w���_��s%(��nj_��ߧ���d)M�/���	��+[�H�B9S�hg���{K�r�%�="�>�N��c*�$��YC��^�����޹�66�V��p-s$y�Jk�bI4;��0,xP��5~�q��r-����=EC��M�����:�6ou���F��j�?���"��ʍ��ҽ�q��&�O�a
`j�e�{�ܤ��؄����f�q݌~
*§�m�A{ ��-��æ
q��M���y��t�6w$�PY��!��k�3�N2�=)�B����,�a��/`�?�z@>�=F�%@��u.�x�|�T�sw�鼊f	��OLX��	��=(�,иOU��E�����;�u��`�c��lw}N�X�v��j�FF'm�՞�A=@�_N����}T���8:���wdn�N�:���y�u�n�ذ�S��A ִgi�#�n����y<��̜�hv��6:3;�]�C��m>�|�c�ݼɯ���.��t��/����,�[uR���P4*�_�)��: D��]J_�J~]��A��e��GYTǰ� U���������5����ԙr��5����u�o�ހE���V:����$�~��M�^���꫕�5�%�5-�5���u�96G (������=����Zf��('�F��|oX�n��{��yZ�l��u�:���j�=���Y�3��x�?��9��Υ��>�~��`����>0��d�O�>�[P7�Q��Ipͻ�m���	���§�O
��4ՎSB�������os�:	v�uʛ�S�x��P��}� V����5����,�T|I�̊e]5+����PO�Ӏ�U!'�������1���Tr����L���fC�EԪ��]z��^���J��h	bǔr��6v6�p��I*�:�n'�G�Ha���o�������'x���_���D�Ї>D�� k�[H�n�nb'}͌����|�/w��v�@�8��i�N��c1�F��.j/tթ��#sW5.A���6e�hd�I�n|�?����N�<��<ڼ���k�u}����K?a�/k돰�������;ȗ+���Rgp�
�DЕ���*#*N����^%�
��h��CD�ե���S�j��(/u;��M�"����o�Ԋ�wΕf�w�׫T���v{&�-%)�,�;]o?=�h� 8��j�qzR��Vs@]c��X��iⓟ�\8u�+k�����X_�E����e\��H-|�]�E�7µ���q��?w�r
o���eLM�b}{�sX���Ĭ�\�\:��P�
�G％ z"6�%�ۦ��['�i�������$)��G�)�)<Z\B,9���4jm���3���Ds�f��l��W_�;W�X���3g��k�p]��{���.�'k�I[ciTK�OU�%��Z�/|�/�Ϧ�ࠁ��ih('�'�8�2"�t/��i�oԅv����Y�Щ4`�2[�mxX`x0�C�j�{\�@��Zo�zu�
(�iE5|�F�ɔ �94c�vl�i����dT�UKu+lR�[��|ڔҖ\	*�lQ�����5�+�)�E�QQJE$/>�����	'�>�T��tjw�`͢:J�<2����,�t�dM��j�VK���=�Nh�ʹ�fG�g��A�w����ND���$.M#���Bn�R�ZѺ���җ��  �wUq�N�����[3�#@'�]$`�w�n�x�^U�����y�Z:�)膡�n,dp��9d�-��2Fb�Z�6��X*Q�F'�V��)��
�(a�$�������͕N��qQM�#F�R���:�y�����K ���d���le�Q=N#��x�A�g��k�ƀ5�5�uuK��5#<O���B�@baR��Q�8����q���=�k>�����V���������A�S�}��nyG/d��-Z�7�JM���/eP�J�(bI�æZW�ɳ(q������c�(� c��c�c5��_�ﴔ���?�G����I� ��t��id(�h,�o�*OA��㉏'��<�N��p�P��5�=���T9���6��0�\�
{Nay�u|�	��
ww}������$v���Ph�q��j<��Q�w�F�P�����R-�h(��j	2����6��
T�116aa�f��P̏�ջ(d�(f�Qʮ���)t�T�c�]8 ��F��!f�����o������<`��!��׿����_G�Ҳ�坷x�L�ѫ���TJ�h�H��1{ ��9��o�G`�=l�2ҫ�������ߥ����t;�4Q��2>���zˏ��Vp����"^88�F_��u����l��G���d������kX�X�3rYjN
U42�>z�^*�:��R�M��(�{��O,*��"1g��hj�=�@��^H���SXFA�x�R���������=qyފ�8�N�@�s!�Hˀ����`$��c��	L�G�����?���*|����Z��\xf/��qLN�C&S1���O�5�3[8}�Ѽx=$	��ۿ�e:!A�WԨ+�����칭�I�u�no5��=�p�"�)n�y� ��� W������h|a&��Zǎ��'�l�h����<+.�J2��������s�Y��[�{���,r;kt�:6��E�Y*�-%&���9�:s�����x��#��[�q�!�}�;�=|7nބ�������π�p0Af0?x?«g���S͞�_�7C�db�6q��M�!��0�Q2`%���� a29<H����	teRiܽws���:��C?g	��,��wyH����,����~,�����t����?ޮ����h���rL�ʸ9��!RtT��J-�y�u%��!�W.���G�%�0��g�N��q�����/��կcTm�[��%�=����-���{����CF���"'O"��hb��Ќ��0��׫X�Sӎ$3�}�@�c3y;��}��Ԭ�u'QNz��9>�	����7P�B(�Z��W�%���C��rʧ&p�z�� e���@}�h����Zw��F� NN���4-�T��˚A�C|$εUm��r���V��u�Jt4�f[5��st��V�W,�p��H��yU���qT���훑�M�R�q�SC��� D<E� Z���:��Z�]�!������\���i�pP/h�p/�h����1(�Ys�~D[�S:A5����f'|F1�����>��SǦ5k��|��?�o�
s�}>�9؃�>�9Un>�������w:����O�'>���$"�r�����q��[M�]n�\f��?�z��vx�:��߿�|�J�Ȝq�u�n�O,�p������v�p��}[����G�|>y�u{q�h��K��TRt��3(.��<Iy"�v��a�G��9����3���j
�XZ��/���
q����T���1*X�RMϿ�MU�����ldE?CC�;X|�a��^���~�4�vjH�11:c�iy�=z�^=r��5v�@�e�z"ᝈ�`{���S4������}˫o�҇B�=l�k5�7o\޹�'L�\#h
��XH��^�?���,|��R;�vOJQw���Y�����ATH��~}��EJن�1*���p<a|p��}�bR�k;9f����$j��2�͖��-B((���)�Rx"V����<d�A�{ N�e�+�"�GE� �Hho�y���@��կ`d$B ������ݝ��6�a��=aӥ�;t`�֨йQz��P�;3sId�i!����K4#�.A�p��+m��D0���Q���	�=�:|��:���:z�.B�A��f���Jl�Zn
}/���
�z͇��Yq5�G2�#�kE�r�:�� �����0�����)��Bt(Fg�f]�8o��6��O�aIpM�[��n<��� l+�g�[s%�}ff��(x� ��E�2F�2>z�J�?�w��e��d�2"@�i�1���8����t,�c��G�:6ŷ��R���(A̎�*�M�������Y���69���ȴ1�͖5�HuT)��7�Z��L�LY[��uE)#g�a�����`%K�{�su;�.T�HQsz�"��Ԋ�*����>�a��gN>G ӱf���(ts�DPoV�L=�h�A`���cp��%�
�|�W�N!���A�v���:_�נ���t���O9Rߩ�/��V�j���QW?<"8�=��\}�992�J�������ç��.��:����sX�R�Bs.d)3�:�ӱ	G������(�r�[�0|`=�w+��>rs���[Nz�Q��7 W�bٲB���:V�(p����A�3�n�5�er�>���qS�v�ݾ��Mߕ )A�@��rԑ�p 1�|��E�:�Q.��B%D]��r+���{~�y�	q:�j�̶�xJ��A�q�J������R�}k�Ä(蠊�S�IćP.U�<���͉W�C�֋��N���UkBq|��p��>��c'�~��zN�>���ʞc��z

�O|<a�q�������5������J5�"}��]$ � ��:���e����{�m2<t��F4F�*Oc"_N*�s�G�l~b#I�u�itq�\G��Ƹ�<�:�!�N�zT&q�5�+L�K����6��QO*�h���������������&(q�p�ڷ�`icq����r��O}
�����Z]]201>1�ѱI�����˿�Ϟ@�����}�﹏������Y\{�>�D����7�ÇǱ�}��v�/�[+Ґ�q��Aܿu��z
É�M�p����~�_!�%������q�edr���H�0����p�*ʕ6���6	ċ��Y�<%S�|��V��%P�Q��N�_�Q�|�kOϵAc$�$Z
}�K#+�)�<��:2i�4�L)4��!ӔEo4��j���ӧ�X-ڍ��-�'С�Oe����t����o
|���W'��������~���^|�<޿~�@�����%�x���矷:�t:���%��/�{���o��_�2<�4Ο���J��7��O�4�Q�n�1i>�}ݩ7,�y���&�9��Vp��c29��7��C��+gЬ�Z�k�D�F���M�����`����h�wx^�l���{h��v���x��E 6cu����7n�p��w�*`�����f��\��o�-2.K�wq��%�{���������ff�O�"A��7J����ӧO�8W�L)V��A�Ւj?X_(��u�:�p�=���E=�y�Y�K20�>�i5:wz�np�{-�+[Duss�&��hh��[���W��g�}nf�qTPז��׽�z�N�Vs/.9ս�Z��z�X�����~���9�w�m6Խ>h�R��~�P�IG�pQO�c���Rw��o�_crj��!K�.m�5:�/?
#L����n�[ŋ�똛B��n{����ҁ��w�u�6�W3�Ua��庩ְ�k6.aO�n���~˜�J�i:&K�562n�=�j���v��K?�|���;��ŷ��G>���˸��K@)��a:��l�@L�Z�v�E�6�����>|���+%�8F�c�lgq��Y���k��95����A]����e��-����ƷA��һV?ɿ�{us�΃_�}��e��e�Z��@Q�˫���&�`1OY#X3�[S�ܻu=,�+j$5�)nu���� � u} ���+W�7�:�����ާ=�!n�;]d��5���z��\����dv����!�ҁ��{�袚y��(�,��]�����f��-<=�O~<q�����6�p�g]��O�\
�� _���9�0�䉩Ø���å<�k���9�.���h�V�o���cV���+�Ècy���w�g�ai7K`Vŉ�i�8���+ti�]>M�
ң��
!����Yƙ���ZX]_5O�ݨlc~�޲K�Ul��Z�Q�Mż�>�'��HV�7]ő 6�9/���[_(죇��.M&��J@=g�o��8gqw�[8tt� ځ�w�#1& z��n`2�kf���P]^�:���"�b��]Ƕ�j[4��ɓ���X���/?ZFj�-�a��.�o�/��G;�4�����bs{�5o��*�����T��K���,^����m��<�~	��R�ɡ���Je�L�q��x����/���gs������K<"7^��������U7�^S�Q�Auh2��Ĉ)׹��T�RQ�nO��^����z��ͮ��6F���9���}�"� n߼ad�3��tR�p�j��m˔�"�/�cfZ��a,�����Fd�?�e9�٦s��h�<��N�&���Ma::l��v���d߇ �[�Fm��޽�L��F�����,�\��a$���qt�3ʯ
6�;��r��2��ǉS/!:^�c{���M'&�*!�]đ����X�N������R�]�Rz)�_�ￃj͏u��C�=��~�L��j+:���Щ�N��Nb�v�6S6�$6��Ӛ	�k��;��^�Q`J�I���7V�6��?[������p@{C���Jf4E΃h�ch(�򘝝�����q����2Eڷ7w��*c��`�M�x��4�N΄"��?�NK��y��W�8��>͍u�������q��1Ш9�_uJ{)�"�o���c0����ݧ�� m��;}��x��;�W���/A�U�&#�$]&��q�K]����{���	�9����4�)��TcY�sD�oQ[Z$�e�I�`��s�<R�;F�"������M�8�	��U��#�O�;������	�	aE�Ռ�҄��q�iZO/4��fyѿ��	�{�-ĺA<w���#�6MEs,�5�l��=���)�2��Ct�������n*G������p���6�6m��F'���(kn��e�5��bSs�5�K�Km���\�^g0�Q�E�<�}c�P�m;��s_ND�5`6�c.��a����ߞ���z����E��ͬ��lX͢�3HG^׀�A
y�VӤ����.d�6��9����W�3�VK&>J����M:1k���$�O�'?����Xqt:mwˊd�G]��t�a��%�*�,b��7�������D�q5K�D�.ceW�C��E�����3	z��-U��v��E]x� jTx	��DC!z�|K�ݲ��Zņu�ml<D�Ǎ�]�}%7�N&�{��i�,��/�@u��^8z۩2��"N�Gd��k7o�o�������2�����D���!�FE�3;2���;ئ�x��@�1�1vT>	�VMc�J8p�8�h����W�p��.�����	,�mS~K���]��~��&���3�=5�<Z���"2�����]�����f=I#�@>��}�+�q+=�a��m�D,ꧧ�1U�&f��;6KV��O#ISL�ШX_�� �r�1��Xto@ӳ�;E���Ee!T���"R2�2��y�>�&�N����-�6�a�;���س�D��R>th�R��U>^z�<�~��޺A�@6��3f��p׫9��z�5\�	��o}��8�� �G�ЩP
Ii�^�7���RV)+���!X<s�Ƈ&ht��lf
���F�w?8�eq���_A&�L�/�iX��Ө��([���=������b|f�x�n}�`f��i��&����'����K��<�;�>�¢��Q��H)�J��=�P�(���z����[�ڟ]Ƴ���-�u�j������9+P������{�zL�,�$ &$��?�X��Ϲ^��w)kM�8�5��������?ɐj%��={���/E+�	T�?�k	�	d���\�	P�Y`�W�<��k����t�u'w,���Q��dU����U��f9�w +��8�\�G4���}o��(Bi���EjPZH�6�z����{�~�Q���w���8x4�I�J%�5rX�@���̄��#��!~R�2]�舂�Zj8 �Pgv�R1�=�+ꥡR��oЁ��7Zt
�1Z�� ���eP�W�-�t�z(>2�%�wV�'ߺ�O�?W(�vY�h!�j.�ύF|V��(]��6�u���|����ǹ3���g]�>��{$E=짞�Z��Nπ����Z�,��~��������u���:9~�w�Np(:2�դ�W,�lߪ�PNJ����3X8v����)?:BQ���i�$;L�iZ�j=���Jf�<=�p�y�~L	�-r�J��u�{�@�R���������${���~W3l���{���Ǎ(�?�����)�J����N<=�Ox<q�P�yQ&��~	�q��� ��$������N_����/�~����?�C\�0���;(�w'0Q�J�ZD8�D2��SM]4il2�ws���w	s��b5�E)UB��,X}J�SAߥt��
���.�3>�#q�:���{u)� �Rp�����聿��O���?7�6�pgq��N$V��A*^G��+[�V�%��\��N�;��[-T��	��/�Ak�A"�����S���'H�clv�Ko�٪��y�ҥ�QŨ�<`HF��=��:g��I��m�����k���&hj�|=��+*N(�/rӞ�i�ц�Ml{ݽ�	A^��2� )��#���=��-�;J#�����"=�cS{�+�|��!�K��e�ed�.]�d^�'�b�4XI����+)|iHe�|>�w�)JkE�E�#�_Eɜ���-_5�H��(h6t��D��`t�w������Ic8����f��v1g5�јb:�xrdfc����;<Ȯ�M���1<=A@8�;�"D����N?���.]��~�
~��y�J�q�T�,����������_��"pNY3�����
4�w�}��>g����=O��Ǳ�9����n��0d�W��8z�y�j�g�O���n�ãV��g+��&
ѷ����1�!��״V6���D�kF%�4����M���@����������tv:������ާ4��X$�W��k��^0�*��Y3�ɓ��5��G弨�D�jTʤSFq��f{��=�r��Kn��՜1��]�p�/_&��0`�J� �5��ge�NߧĉP�K�����eʫ��k p�z�F���mTK�x����180�,�Z
6�p�{`jr¾� �� �kP���#�O`P���I/��9��V��WQ� Mx�H�����.2�<\�Av�Nu���1��a��]��l.��7�ųgPl��E(�]x^K��mQ����&ez��gr+�m��'A\�����@�W�_�aǠ�#�C�lX�i�EpM�Hj�"�'�Tbx�Z�N�iL��#���^(�a�7r�Mm�KG/�3�~ɱcHo�$��~�.$�Դx�SX#d��u�^�sZT�3��jխ>YvL�X�h����Bj{��5瀈Z�ZP> �,q��o�?���y��>���y4Z��F�c��t;>�Z��uK�Av������*��>=���'�C0�k^�^UG��*W�UC�&��������� ky�=*�u����&�Gl&q�����)�� �U��vC���rS� zo��!)e�mF|�����C:WF(|�vx<�ULO�Tm���g1wx
w�ݳ�|å�>��5���6^{����7W,z"���{jf��ec��C���ɿ��Gi$\(72���!@�!�������x�9\x��^���ǿ����P]1�Z�I�ڴgx��,24�x�:f��3�(����7��tf��	��# P���|7��{{D��B$>�V�m�7�l��L�(R���N�w�c���V����ͩVa���7,�ݣ������� ��%�^�~����k[�k�T�?�j�e������n
W��k�$�Gʏ���D�E$��A�g4YQ�A�*i�&�(�X5��ad3;4�C�L�L�sQ{`ry�����t�+m������\�&һ�U% .��PV�ņ��Z��c�`$G9�d�h�d�5{��,1�ҫ�����k�Fb����γ���8v�E�����
��˔��n�����)���#2��{�q��X۸k�ܥۗ�d�q�s�w�xp�!�9>j%�zgO/`3���TcGp��Tip�A�V� ��2�=�F�M9ڱhE��]�}��@�H�3�� ��\�g���>��@���p��9��># ��~t��Z٬���ǽ�Y�Zw�OƆ)j�G��R�������9uh<������s��IB!��;�͙#b���� ցs{��u��o�=萼�{
�il�dO`W�%�L��X�H�ٯ%���8�G��# �Ԟ*e�����Cx�u	�~
!g	�Fm:n��K�y���6U'�as�l]��МQ���-a|b^����)�;�C^��(ZR�j�s_�F�@.[A���LE�'�`x��?��sx���P�+��� �gO��W�;X8z�R��`�o(Գ�p�&p+�f{�ϩo#�6�V#(�E�����1�q)si-�����Cݽ���n�5��������VޜӝME���?u��y��[���b�����!��L����O/�WO�X'��4"S�1�n�k�L1���\s�k�笽�C���L���p쥙��+���I�������p?zh��g�yLEc�)���B;� �>~}θ���j�k6��z�)%��㉏'����A�t
�s�C%Gʢ,�C�A��!���ױ��:������;�<  #����S�|����ˁ�J��<��8��#�f�a��4��2["����Q��( ��B�$A��c�IN,��k�0�WX0H�WT��>�S?�L9��l�iX�����=0��G+B�T�������?���5�������җ�>�k�������#�S���!DhL���7��!�����lc���C����G�yW��� 9r�@��Gi4���xn���^?����oݢ1��'4�@x�csT۸��U��L� M���Qtz	<�������	&���H�^n�k���C���e�h`#�Q�Oacc���m�e�0��4�������{{<\�'�Z7��۠��c�fRVx�=+���MRThey͢�J�Y���˸+�(��H��(r��5�D Y���S�YS+��Q
^��|TZ��S�N��G��?�y�]l�OOL��[7�BӃC��ձ�p ��~�?�"��C#���֝�03;oߍ�[$�N��S�R��{�$i�]������Ҕ��]]�}���;k�@�� �F>�_��"�	"	�� W$AX�.��3�czf��������*��:����@A����lwWe����{Ͻ߽�̌O��f)c��i��LU�5b1t��-�}����dB89{��1�L]d ����C���O87�4�Yd�4�y�<!^Å�g.a01�y�>�l?����|��އ���H�8�j�C�Cl�]���h�N�����Nadb���ҥ^�zR����x��������V=Vh������*\�ҹ({'g.P&���kmK�A���a���.��惲wʪ	hhkX@O�CM#]�<s� �����8�Ɯwgݟ����g�m�)��9*�[ҙ�7����~���yV{�j5^��;;�Ol��[����Loxp�@�>m%����O>�_��8��e��I���~�l�/��ս҆��7�����g.2��C_��N�.n��o8�ch������3P͂s<L��1��1�ŭ��(Z'}�׍���Y��]����8��l���K0[���G��Z�Kzoc���$�M�w��˘��<��x�d|	��d����#�������Ռ�{�˵�,"�Ρ��!ƣ����"�������)��x��<F��ùӧp�Q�{�@�d�0!�)�Nkz��{�}��K�i3�L�G�E}��\�RGZ��G���7P�{����2�9�8��2����+R�O�x���MEH�C��ү�T��}��&}E���s�)Xu��툌��d�W�������Gۻ�Nv���G�(���C@��8�O�٭5츎(j`~�P�M' �<���v~\2Q��Z���SP������\�r�1���8kt0����B51�s�z6�h��QF����ۋP\��.FÌ�\qbȀ�M{�+<n3"�^�N��Dȍ0�G�nI'���N���a��J��?d�j��F��D��]�/��Ob� �>��Ro/��_G8N@���9��d��`��9i�u���V6�Q���)���S3�����x�������ş�%�
������x#_�y���p.,J�+�����c?���폱���W�� ���(\���ays� �����`��̓o|�琜����>������?��2#�_0�׍�5ܝ�k�ٗ~��a��U:�Rs���/��`k�p�+��[2�FePR�~��!s��"���fu�F:���gb^�B޴���� ���K��������"Y>��Aƺ�,�$ �'CW�6�'�X�e�e�$?91mY����m��>�<��zäɜFڶ���2��'�������`��`S���]�����}�.?�R���!����j�<w���o�ƀ��f)��/������"H�Z�����cēQ��Mс�b�(c���A>��aln�$"8?{D���H&�V/;5D����,3 y��@��cY�CN��J<*���
��m�8&�P��[��A{Hz�H�������W�� �q�+6-{��%@@;12�t��p�c<�rÍ�S�����Y�2BQ���n�N��N�t�����Dέ+a���	��T@E���:ǽ�w�ߺ�5��\��_�����tu-��I�����u����S}	��@��Tb��8<���t3�jpR�Zח��郫V2�9��g#���m��V�6q7+*0� F�,`+�{��}\�z<<�~�9[�|n�W�X���kJG�r;K۶�;sb/_��ȵ7������p�r< ���������$$A��
��Z��s(OG���"�s��-�<n<Z߄��w*>�j��%�t�т�(Jg�����h�zƍ�����8Br�H�`����&L=�R-����\���E49���S��'�섣F�<�?��-�[��4ҘJ��ҏh̚!�8&'Nbqy�+V�=I�*N� �������ö  ��IDATmģ>n��v�@/"Dݗ��V��B���Պ?5t3py�:�zH�4�5Ο����"gƱ�i��2�j�
�D�^T>�j8���9�ٓ�H��hD�m ��XAA����S���6���$��fvt3����C�D��(� E@v�_v}�b6���n�P�XW����r,��r�)(|z|����ܮ�[4!m's�]h��U���jC\]�����n�AF���x��3�=�5��@8`�Ң�r��sx����c�^�ڒ1��G@R�D����V���V��u�ҹ�<�\��4�}���˸wwI鱺 �2���}���t��yLx����=5�g�^�/��Ϛ����[��7��u���."��C����<���F��v��2��&�����P,��c���6�c�����`I�#�XY������3r���p��W���K�:��U��K��G@�S�%����^�EP؇l�M 3�kϟ���5��'����5
�{���R"@1mL�^>��h�Q4h/;�N$0V��q��n)��z��6ߧ�!OUV��][��C��̞��7;��' 'g-'쥃]���^_��}��v�{�y*�����N2���ZLF� ��p_��7m���~���tΩ*�� Ο��0�O��'C�QA��F�Ǐb5f���=���� f�O��fP���L���!��⫔q��C��
0�	��ON����W;淂�� �����!�kV�|�V��nK�c�(�n�����X;X�w��Vְ�t��	�s�V�7����o�zUO���;�t��$��0)���;�?�,�.?����Ķ�2��՚�A�X�����)�t����®ܛ��2qr]-W9Cm�v	�E%# ���6��S=��X�g�}fsId�jXQSQ���Zk=ٲ�yfc�ֹܥ���ܱ�|ת�#�YGVtDp5�>w��HsE�Hݗ��͛7M�L UY��V��1��_0|D���L�^-kض��Ӏ�����d��q&����uƧg�&8�5��?��?��_{��w}�~��=�KW����R���c4�
��c�A`���3�D�S�)��X���ky��K}�~"R@)_��-�t�hi��Ј_�@"��&�Ճ��������1�$(nx��8&��q����x����1=��D� ��4�=A����M��<�/���P��66v��8�
�@<��+���;�0PO�� ��5 ��r_�ʀ��A����~7�R1+
{��|�c09:E��6$�Q츬�N[����.��1 (m�=r���G�؉�"v�Z՘
��,���No1dt�m�d\*Q��v��6�=NcJ��в��1�sj��|� �'
ɖZ<�Z}ᑿ<jL1 �8l[	���?_���l�J������?�z��m��uђ4���8s� ������p|!PX(�]�J��$P��GB�^sb!�6K����
Ґ�8Q	ʂNM���n�H۔ќ����G4���p��9����A)�VG559��%j:��?�A�A'�o��� H�Bj6�&Q�a���#L�{�׊�!�9��������e;v� *G'O�]~�I�x	/_�`�Zo��usNZ�R.x��7��Y^yd��>��cx,�Pl��&%�T/�6������4��p����_��8a+��$�A1m����������_C���o��#���SH�`����ML� ��`is	��}#�v��LǪ�墜E��1+�W���Ei��@E��b�ѺS#�����Z�B�*ȗ��eG8^�g�3��+�	F $1�X�W�0)S$�$�&nD9W�u�ڴ����@�-W�G�[Y���=�Ca���2唝�<�ҵsz,k����1����O����;[��?7vwvP*�0�������i߻�҇XY������/��Dw?�#�pe��k��@XE���m�[��x�a;��p���ڃ��!΍�҉#��؊X�`?�59��#�V�.j�����*s~�600<j��*u��M������ǆ����{�ch��eʕ<��>c�(˧LNO��<��fz�L�p�G	C�������{8}�V�P/{��,n/AQD��Gz������z����Z7xր���֙��tu�p]�
N6�e�JZ�����_��l�195kپ�h/?3bY�Օuljh�Z�pbj�怶�'&��s����6fNL��g��bu��F�T�r�`�	"6����X���7��pX#_� �mCo©u��>n�A��6�h{Zv�X�#���'�i�|&���`���w�r��p��)����M��K��x��5��������${�Q��v�����q�-q��T$��k&����q_]ZBj��y�r�X���T2rw�}�6v7�hu�X���/^x��~M`��U�/>@�`�#)ܽ5O[ȵ�D;P���W0?���a�|���O>����S��3�ۯbt�$���[�>�an�ό�\�_kq}m��vrW�pjz
[����m�Kf҃'�Z9��ܝ�B��6ucom�sUD�9����
���pL�wZ��^��~��U���\��4.�������&�P���Qk��t��Z�B�� �Q�ת2���5����em�Q�p�Iױ��Vgo ��j�t@T��#���2"�+Ie;G�ѹU���%7�ֽ�t;p��dq���uˑn~�i����/
c���3��	ڄ����|� j��#�4/AC����I� x4���+���E�ѭ:��>����*hT	�pK�Q����ԩ![���h��F.6HE�U+ >�����gU�_E˕DO����.� ��Av��ϿFC��\}�&���Kw	ؚ��ߙ�&A��=�����Jx����)}�[�c�Cȶh�汾����&&�x��bă��>@��M\��2���u�����5I���-LMri0ڧ3���3��}h�=��{������>BH�a}��N�� pKc^���c�!��+����]�t����w
K���{{�'#a�������AK���LȽQ���]ۍ2h��Sd,@(c��9�#>�f���7��FP��{ �;���DŢv�104��C��x`h����#r�����[*��1-�Q��Ge� E@���>���~����������\K?6����]�[_���>�̬$	������`p?�gQ����Q���7舛�K�L?[Ym�f��9�Q&���-$8NM�Ӏ��������A���(n��y?���d�� шU��Rq����ܮ#���{[��@�X���������eUW�wP&�D�������Ex��b��߲~mwK_���d�cܓy:���9��*WV��/-�P�φR�6��bU�]uN��~lם�;��9�l+k���9�5�ol��'��!:�R�h����Y�rVÉ
��F'pb��k�O���^��(��l�c��P�[@Q�L�X�U�����3h��)Y^^0����ވ���}���s+�PVS���(ŉ������G�p���8{�,����w� 1�J�<W��`t���0q��z15~M����9���
E�\��H�b�������~��G�`8Y��q��\��_�+�C������B*F{x��D�����79M`�����i�����$���_�5���>/�d�fWc��\��:"�=\��½������҉�@}�X�ӯ��S���^����!�~��I�4�iK��\;�qrf��R�4�(��l�EG
%�:�~S�Z�[������}�O/�1�����)��h�>N�~箽oO�v3�������� V>��'�<��ƎH��hp|���V�C}�fN^�}]G9��2�i��D(�5[J�7� �ܴ���.�K@5d��w�#R�0��ˠa�����j�!W��为�(cZ���(t9�u��-m����܆/�7��6�Dd��w���I�=0Iϸ�2{)Z#���i3n?��X��7�r�g�0_�i����>qA�\O2�5�Ԫ~����ߋ~z<=��/
ۑJ��K�KT��h��U�&�BFJu�h���ɜY��&�˲�1������	�"+�˶u%��B��@D\]��hI�RYy������$��Y���W�$F�=�*{�����" ���pv��s�T]&��᣻Fq���Ψs��H��1�Í�?���?���"#��cN����o��T��m<�j�ӏ~�WJ��.���.^z{���~�&���7�F�}�gi���;61��]W��h
���Q�6�/�p���÷?BﰑJ���KG���n\e�<�߼��.`dx²9k;ydKa����m=���!�ol� �V�N�����?�fxD͠�Q�x�)��C����	0�Iw�2��nH`Mz����w�:4S��;\����2���܃y۾T�QY�n���~�g�u�h�P��� �z�MSZ���M�泏�k�_��FF	V���79��-����3�����M�S��p���H�J2�j[�~:Mɗ=��X�K��?8ıڧ��KϽ�<u��F�F����%��l�,�\���ci>O�-��?y�Y/N�<wC]�+���=�b�σ�ZCIu�/ �u��нL���u�
�^}�G��(��tX��ʕ������k�gN_ĝ{��d�\j��m]i��R�'���z�ZO�5�|�jc�k$�)+�����Cv-'��]�0k�y����-��̚v�>+Rje&Ug�9p��m��T�Q�׻x�.,�n�&ח2�a��^cuyՔYt��C�
Ҕ��}�A�^@MW���Es�K�+�57����U�&�%}F�K�k��C��(p�`���mFGeu��swm{RM;��-U�G�>���)d֗M�RM]�:'����(���8�1>5��D��� 09=�����m	񺙍%l,�� f��8J�X��[�{��|�8����\C":���"<�6p���^����h�6��b}�{�jc/�}��>�.�y�8l2�b�1�����87;B�ܤM)c���_��g�ft^�@?񵯢�����ηCDCA���q|��u@���cz|�vA�G�?�\G8��9�&��>	bnd��n�����=R+� �md�� X�ǣ��9��_zÒg=���T��Lr�V˴SA�pvu\F�I4ZR�5�
�{-�(Bo��3a^d�w����'�5.�mU���V� "�����7Ri�O���ǚXԬ����8[s���vH�;	-T���2����l5��CP�5��)�(K("n˓l�֨��~�u���K_���KS�F@m�B��.��u��19�hQ-׍�$H`R�4��F^:��:۪}�'��t|V�!�Ά�9M+�%:0���m{�^�.��ȥ����٥\v�J{E̞C�vL�h�-:��8vl �{��H|X�_���*�g�4��i$C^�/�H�p��I�VÃ22�>?�_����%<����7>�H_���J��6vyoEjF�P�y�f���_D��~u e@�F0�ϔq|h�A����{�ࡇ��m���QF�y˂ML��y�1z,bzgs�caT�e:��b`0I0F��A�J'���� r�L�N����1t��1�stu���vNБ��R��Ϯ�m���u);�uX�g�~&��h;�]��B6g[�t&�	���`��( 1{�S���1�<�ݳ,D�����έ����6�	E�LL���c�,>as%��F���$����]�ޛ��t��b{cٺ�CC&ť�7�É�������SJ���;I��py�KK��4�y���$��?�����
>�h�>�-�s�q���}�6��r��n<X����%|������1|��A�$�W��Q��_��H�FQ�`jxO	}!S����?�A��G�݇��א�� ��
��h��~�m��z"Д�N��e��5�E?�w��VS9j:�ѡ��������MG�G_�1���jG�֐14�l-�i~�WM���W]=��X���c������(�ۦi���nu��\�n�Ƴ'N�b��Z�S�P՜S��2�}}�Ƨ;�l�3��U����/賚���q,,,wb��@� �dޛ�G�@sQkBr��:�H&�D,n�2%-Y��d�����|p�x/�{7����ZM!���6����&�{�]��ck=�_��_��Y���� Od<ۜ[I��؉	9��pս�0ꭇp�ajH�eY7�&bIڣ"���׋��TC61~������Bh�x����We:�1-dZVJ�+nr���fi�";�Sg�"_j�8��1=t�A�9�_���w����+k�p�}A�k/�r}�ǐ�E�PC$A��c���^�>� ��!<w�q�*%{Ʊ�8�آ�Iq�E��DP�G�V-Z�i���"�UI@0l�TbI��նʎ"F�]�3�ۢ�B(8��c�T�
��VP)k�0�hi��g[��ڞ,Q�K[��ZǴ�E��@��V�m�����y,��D�)�Z�x�����d{,Y"��qD�meuK[��Od�p���fM2�ɶu�v���?x���O����A!�S[�j����^���ۨTcg���"5�tX���tLmm���v���	U+-���`S�<���{:V��k[(��T/�X�M+W����Չ����{b�0����(��"[�=��$�S��4m���4xO���O�w���m�kh���/�"i�FG�f����AI2���rKЈ����99�j�d�)�h��y^/oU/�Z$я�a�`-���������`ۡͪ�R���VW0:<�h0�����D�8w0���Ĭ�$l���wQ��`��	�[�-�{���9��Nˑ��f��]wO� ������H�G���u����BNU�®Ƭu�Y�����}v;X�9S��	�3���yVW��v�����3�|�k@	��c��D�cH���eck�j�"QE�9�85mt6��mL��|TsJ?���DzL�W[u���D��6]N�~��cl�N sIu�j|"��t�֗~���!,=~����-e���#{�����m�$��i|"Bg����5�x�ny���ǲ�j�|��]:���f�>~����ӓϡUhY�e��q/O ��O� ���$�p�j	?��;V�/���R��茀�c�w�:<�EW�A���ɓ������X��K0��Xl?� �<1��l��ź�Z�l6���D8G�}�:Yə�jH��j ��p�ݰ�[4;��A<z�hTER����T�@]��C�(Т��@��hh4��ԜrH��1���}Hf�<�bŲ���2�����B��[�8����,�^5�/���׾��ap|hl����P?Ay ��!mU�e��\�/!L���א�}��vv� �����g�-�����ݍ=��i+�����1�-���y�����t�8_�+��>Д�de���`� ;���!��1�8y����>��(�u5z�	��^vV����lX�%������7$�+ uzA/�a�j�	���+���Ae�XEz/`���h�-�NF�uGm4:U�d�8��^��4j�
���XzX����o"�څ��E2�{u���z;6���"Au�;��\
�k�\y7Z�����._I!��1hX�I�alY�p�}T���� �Sw��%��L���������ێW��*��r�a|���ٖ������x���n�Gm7��|^�HyE�O���������/u|!P�.��4�q�I��
r�?�4�jb-�W[�j�(�D���^A�(tn��8vv3�e�;��.�궘%,���դ�y�FͶ���,�$xt[3B�Ƣ`E�rB�z˜�2|�\�������	�[4 	:�"��F������qޯ����4B�H�t����J�6g*&.�ٙ�y���~���C*���]o��될�N8�w�g�<C�QDԗ��h���ӏ��6���2����Va����O���Rb?�gya������n=t*zW����c�����Q% �86��]�>#�n�t�&#������&S|�3��)�j�����?'��Ӝ_��z���g�m;�hXY}V�W�Bן]P���r��\�5ۖ5��}
&��:��}Lu�.XԶ�>�nj?��GKHy΅ �A�ɛf@̞:���	:��쳏1��r�RX��O������ �P�5��Z�j�s.��?��s����ɡ���p[9��>:�j�2�ɩ������&�iqeN\$008��m�;d�1?wo�󧜃i�'��=����X�O003H�Q" �A��E����vnN�&��������F��������?2oW��PС��ҁ�C�,��#�����mtI�m+��|BG�f���j gf��9�W��Wd��jU0h�֩��He�D1��������:��I�d�nlo8��� [�T��|UKi;B��\�|��4k P�׺wQ����d#N��c��e�Z�O�jF�"�5�����|g��W��uVd�,�ΟNg�;~����3�oM��4L��i��캱8�>B�;�Bd��7�|��V��k��ɜ�(ꝏ;n\�>>�d4w�]�sq^�>�޾8��pN�WF���i�����L���x�wP�����x?r��r8V��������Sp�9ݣg`�G�試p`�.\�<g�c�C:��h���K�?�|ˇJ8�F��^WLuW=?�|/����ɹ�C`õ����zi��s9�Цe9W��\���&��qfz =	J������A�v���\'x�ϴ��xc� mo)��F�ɠ)�W*;�������`�5��	h��?��1?7���Mw�_Cӳ�t^�a��f��!���:�5�8�;��s�!���XJ D�>�]����]�M�?w��>V�ްn�5�h[Y=$�N�����*W�X,����4Zm�*�UM�Ӓ���Q�����9�y5�Zo{ZG�H�8��nq��LEת[*���	�.e�g`p�"%꾾����Gz�m,J���F�1���
�V��7�O��&Cє� �����h"�]e�|x���[�X��\lN=��#�>���<�*�R����~�K��=x��Ɖ��e��h���b�m��9�hX�]8U�H�{���٪ȡg�v���?z�Dd}�$>��.�\�4%��,�Qv�=���C�%�x��K������^x�*�.��Ý���]�:#�".^<�h�����g��4���M��W��n�`� \Tz�괮���lj7��l]f�@�e�x��Z?�_��R�ġq�9j�m������f�]��"u���0Z&�Px�}	�v9[9}I����������`W��3��M,?���wn .bh����*����J�8{�9�s����m��9���ʅF��k��c��N��ߋ3'g��	������q���n3zWB�&��:���ɏn8��2N�����:E���Ocg�Np� ���t�A<^Z���6�67�>"�E��v�}-W�o� Y��!Aa��Ζs�s}���H��D���C'v��C8u
�o�o�i8h��G�bl|����}��6��'�_c&P�q쪐�IGu{����r�O�q�/M��S ��3�K�����M;�>���C�?R�����76v�ZgϜ�No9�MmI3X��A+=Q6�x�y�h��h��%'P��7�8{{S6_4W�<�ݟ:�H�<C����=�7����Zw��=zd�\���U�S ��������Dz�{�������y]w˫u�n<�H0ù�b(�%%0�61<0f����%��޴�X���ݽ��Ά�����h���c"��檕�h�\�%���9=�H%�p{���a��>���Uv��0�CS:5{���Kh��h�����?���~��L��o`s���!@�����j(ԶO鹇��r��� "��Xz�����TZY64�5����1,�H�08?݇,�䵍d9g�-�_��Õ��8�Չ�U���9%x�5�O�(a=MZx	���n<����*�#�V��Q.��@c.[�.�p(���(Ƞ�Ui���"6v9wP��=���F����a^��k�bu���$�`[�0��r���`?���6nc� ���S����)&�������[G�?���#@�25�&��"�i	a�Aّ}��啅�4T�޶�y������_���§�_��B����Z���u�Pd��B��\DV�@�(�$��N�F:�"0i��`�I���#C�A���nE�Z`^w�D���gA��٢ϔj�a+nW7���
\8�N���Ƅ�W?W�a� �'�јGQ%�덍ai!�_�ş��_�:�������������W�aB��P7~��:/��-;~��mrh#c�J�!A� &���~��җp��e���O�/��o��{'�������~��5�������h7�^�^���546�����$'�+��/3����0��������"~�W���������ZF�Q���g�6���8��ٯ��7�������]F��C����֛�����կH�X�\`P�^�ޣ��@�@�����������ƈ�Ȱ���d�<u�����q��2���v7S(@"P��:������h+S�*���o�8�6�p��?�G��h�5���y�&po	�~�'��s�P�(���T?�&�?�s׮r����s_��o�>.??�vU����<��`c3�qN�S��R���D_�ƻ�J5��l���Jo���x�*z(U��p�9�8y�s���a��&�lɋ������{��:D"9��c�2惏�+_���������oⓏ��o�d`�c~vs�!��!s��`��j+,�On#�� ��(zS�&����{H0��T�6��5��=�#;��V/a{���=~b�I�{]� {�6V��֭�6�#�c�jq��IW������"�\������\��i���W^��e�Cݗ�Ż�(�2�Zך��G81����\7;���b�55=a�.�{��?�"W	�ȹ��i-��o����Z�B��ϤTŅ3�Ht3�z��D�dݴ��dkA�{����s����CD	�ǦG�ng��_��F��x#�_A:Wǽ�������e�L�6=�zE�4T�L[k��9���g��N��>�(�Fy�խ�<���߻i>��v���G�T#Z�N�]#��`�kɫZ�c�cb@t�@�Xvt�[նl�P3�WЪG�Qc�ty[U��\�4�� .�����BSS8w�uT��+m�ǀ��ky�� �;4B�!�Q\6�!�������?@�p���d�Wė^�wa���w��=�r�j	Q�u��6��&�E�ע�vl�����'p�4����K��3dtr�<����s.������,��N�C)�ut�;\�h:]&��S�V���O�a^'_��C�-�}'��7*�
z�d�|�*�vB\' ׽Y�I��4R��m��m=2�9�`RM�f3M��c0�T׳9��Q#����t~��r��ӆ���:�8y�KIB�W�1�����y5qU�.��A���E�1�``V8[̥����2v}�d�{4��H"w�GO����1Rd-:+cly��C�RrRb�wy��	f�2.��!�1�� *�:1.1�E������0�����.|xcgN_B�T�ɾ!�p���WB��x��Sۨ->D"a�uh`B{	�K�`t>��O�������a�9��0��3��Z��N�e�)��#�ce�>��L�`d���������E�4\�[|wC�J�R([6ś� W������Q�1ɽp\\���@�U����E@�2�F�e�n;��D�SFFY"m�
(
8t�I���]�}����)�'G�C٦n��3��.}�揳��x��"�ޕX��#N3B�h��P]_[Cz��?�E|v�SL�NX룇�����8F#�8b����W/�y�X^^��>��w�/�̉3���p��p|zk�cv��&�����.X�k�Q��u�d�����t�MQ%��"a�HR+{��7}�}y��˸}�1�� ����o�o�k[[��[7~�c�C�����:^z�5��ҋ�X�2���F+��{��x<�ss��l[�9�	�2/��U��������GkD�ED�����J"T��{��P�y��G�M�(wԍ�����:S��ҔE�V���d�v�vS�F��:��l�Lu��5�j�2��/����ÃG�e���ܹ�4"��	��G��t�UM�x"fM�y�Q:��y����{�]K��Lw����njz��x��a<���:�2��r�2h`2���Z=	��U���i�*��e��n�·�E���X����|D�U����g �8��6z�RHӮ|��G��o��տNNM���h�<���6w���C[�u<V���}y�m4�����G;���/��ؘ%Fq�����3�仌�E#4O
A��p�k�J{Y�F��k�? �_�r�����qTNN�C,]�R��`�?a���JK;��SV��;D�`ht`�J3��>|�C�̜��v�W��ᱳ&{:�sO3��6�����P؝�h	�Q�qi{��i����ж�P+�P)���*OaW��'�gqth�scߘ-��-��P����~�|���'�F�9 X������m�1n]q�6k5�k��>�$v�(�0ktZ�,"J.���{*1b�L���5�e%A/�Ֆ�ji7LsQ@�i��8�v<{�(���H�bͩ�տ�6�^.�s���!�rj�#Q^����Q�������/�}̐XFP�q�^6^�z�I�K��X�X&b`��%~�+k�=��(2����>X���O,��?,�{tz	(���5:\`A�[��|���1�1w���l�I�P�"-�T�u˂�0�������"ȅ/]�r�i]��JK�w�r�0�7�{\t��$
���O���9���!�v�0=5�_zo����c���ʙ��Fg>�g�j����d���T?Aj��: ���^�#��Йӹ�96w�4�~<�����&�Oatx��[�����nZ�V���_���Z]�j�j�"�?���)u�n`k��"uݕ+�`==2�����v��e�d���s9�.삄�҅��r�Ӵr���qYS@٢ۊ�'#(�T=jpQ¾��m�L�j{P;OG�Qs�n3is�ݭg�u��K@Q5��>��/���mq>�9&#����������]���FG'�Üұ����|��p�����u�����[�Z���2XA��3��2A����MT[�S�|庈���R���W����pW��/F� epr ޽�Xb:��w�[C@o,�P$��܁e�T7�T�z����>�P����WZ����x���fl__~w�#�Ì*��o �?��L�{�[{�F{1�@'[L[%��[A��UNG�Y?�|P�Vc�-X�l��[�F����[cJ78�֭ ���ɳ��#�����5�|��5�S5��=w��]c�C��uL"�cm\�45:H5����,����Ȯ{{�5�$�(���6�2i�Wr�:]�z&�[�j�vd۶�,p*'�L�qx��M�5�ѱa����u`��f��=~T��xm�#%s�/]�/�M���[@$�[}V���$�1�-����)4;M�Ñ KD����&��z��-�r�G;����eĢ���y��ȥ�v;nT8�V��m��pq�20lL�Y��0���bys��w�X�8U�ڣE��c�4�X|4���o��\קO?�_�	�Ik2�q�S|��;�O�W,lay~�?wcj| 'f�p�t/���?�}�ߠX�B�;3�W���l_|��Z�p���s��D2b5���ۚs�*߽��D�]�Nv�s��*����*/�G��Do���	rԨ��nخ���z@Ia�]1D�;{|۪f������=����/�;W�R�-eԻ��NM�v�<��Q}+�� ����(R�*"a}Pƚ�$� &�&���{Vc_�T�CQ�{l[���"�<'�r�nW�l��q���ֱ��}��^�V��j�x��p�߯���xz�_v:J7�;�}B[�d�hEQS[L�0���%���0#b�CF>՘e]K�4�Q�F���'w�����7��z��x�_��u^�0TF7���ӊE{	�xM՟�-��x��%��VS��O���Ms��m0¥a�e�a෸���s)�S}غ����9}�Yb�8>��c#]Qv�ܲ�q�2e�D-����~~Wj	�hT�A��(9(+'�u��-�����,3x��H����##�����V��ŮkW:U���C\ű��i.��~�o%P�Q��^:��H
-F�M:���ɿ@�F�[���X�.W��01~̊����i�b�Бk%��j�	 ��[�rױ;��d��sG��i&�����y�꿮2�Ϋ�t� ��~y�O�Z,*>�����i���s��}���[�yݍ���٭�<��t���M�0@@�������o�1�pah�>�����7���w��'���t������!@����@(F���c�+�X/�=ad���d��&�ߨ.4tH��\�e������^΅U,=^q��A'N�!�񇹇�0$0�!�����#�%��.:(�j(�zr�_���2g�iWx�C���W�7���f��0��^��&������Y�O��1E���"?��$��m��9��]J>�<����>��(	99_�
jd���1�m2�n��3�9���*��sssFG�];Ң��ݰf.e����Vd_+;5��V��DMj^߈e��&ǘ�y���o[V��5s��F��q���G�T�`�$5�A�sj�Hr�H�M�y�����QgՍRG�o�s� T�<�n?��i��ZKs�[����P�԰�|��"w7-�l�/<n�+�d[k���ݭ�=B$Gl��i.���I����`�վJ���k+�v� %{�}�&N_z|Fe�wvW0П�}�q����'��8�2mN"9�@��R+����9Wv8ߧMF0O!�`lkm�A� �g(jk^�µ�.6��@">��Ͽ�ݵM|�O��@�e*4���)�����x��9�`��7���S����m������/T�cw{���V�{9���|W"�m%������<�C��.d
2�l�_QO��d?k��"߆u�ా�����6�`��6NLY �`rM��ۅǚU�JK�%��zqj��HѤZ.qN�X�`%~q#Җ�
|oEDi� ��6�m5c��u�j
Eo��L�ñi�[Fү��f;�g���u��>#��=��qs��O3�O����@a$�k��j#�l|�����|���y��P�y��!� ������'������/a��M|��s�t�Y����M�x.�"�삊l
�L�����,K`ƭh�� X%�����k�6�`�k����4����g��:mCA��ܽe�7�;Y:�^�?����܊�ז����U�*.d�aܿ7��/���CL�=�^� �8!�C>M�Å}��$k�om/�)Y�߅MF���,���h�4L@e:(�>��>.����x���驓pWi�#����a�����n����$#�������N��UvA���i`UǙ��/�p2[[� � O5}r�ݮ�.�G����ʭڜ���K����8�F��������䙺�Ji/w�l�?p1�a�<��S�|_?1=>������}�����L��%�衃�_�t"�1<ԇp��T����ǀ�3����[p�K8yl�ѐ;t��=��8�wV�]R�?n<��rպҥ&��L��׉�	�Z����>F��g�_��+�Q����	D���Ur���"ǥԃI����!��;��b��m�f��F'R�ө�{�74����5k�UD������C�Kk�<�f5�3�_���)x��(�k�,�/���4zzÜg���1�뎷@��C��iNh��`�qPY�ƥ�4��W�(�Dt]{�}�l��i��~��m+ۨ.e-e�yF;K�g��Fm[M�:�w��*�Y��$x�T��@��E�� �߱����R���Q%�	ac�!��cmm�c����,A����Do� �j���]�;��zO&�� F\w����I����G7�SV�.>7�
���m�y2�?���f�@��, ڣZ2��
�~�CD{���ˀ�s���:U3ki�,����N��i�Kq��[ZD�o��V��tw � S�# )�R����`z�$r������F�a�<B`s������idi�c����N��g5�9����c#F{0�s/^�?��o!e5�b���׾���$��C,�<d ����$���B�>�3g���ƕb�jkY�w�'b3`R=�[������j�8׸Vr�{hp�Dz�&)e��?P��X,;NK,�p:umX�"��^ך�:�-��ɪ:�>g�K�+�L)dY?��s�]�2��z�`�>٢#��j��ѧtZN�q�*��9���8A�d�,?��:Ϋ\_�[ͥ�D�<�h�֚򐔦xNGL��H���������f
#5}(&	e�n�-����bV-.4���V�����������W�x���^ƅC���L�>�t�;��U%PoU��¨1��V��Ek`��,E_��^��%��ϗ*���v�
4���&�V�!�7B@�k�"�S�ؽ�P;EGt,9�Ǐqlv�����"b�)[���C�U��p2�s�082M��C�G0B`S(Y1t�^�+�6i���CF�q��2�
�Ij:�F���V�x�V�4,UD7�v��Bn+�ѡv��l�#ۆrgx�>F�}�!��f�8&`����Ձ�@����հU����@�[h��w�r� R�~'`i�*�'�S6�Kg#�`��.ד�9�j�b��ﻲjv��n��E�t��y���ix���i�=X_ݰ����V��b{s���}A:	����87R��)�<Z�A����o��}Vq��2xH�D���TN���c��_�NF""�SǑɕ,S]*87~�e�v9�\�0�G��P�C�{�9�"�m:�|ƀb��tlC�#:IDJK��h����M��T\���U�;e�<F���j��,��CL|�5Ɠ����N�L�pw��4�&uC�������_���}��;��' P�W6P� �>����K�2.=Q���db��T6���t�7q��y|��{�<63mY@���'5�r�z�}�R�!P0�#u�[w2��gС�*БSU�����M�U?ҟ��Ùx�ؔ9a�W5���>VV�6p�R��j;Z6�5)���*s���~�p�h�ߺg��w���A'����L`g+c�20�AHm�rq�*?�5��� �N8LoX�q�����%xx?�}1��=#aO���$`�Jz5�H�ĭ������zh�%D�Qe�N�����;F�5<x�v�&�hC�Ƴ�zF�P�'�L6m�je�����`�����c3�>��n����������<�S��w��U�no���]ܻ;ϧ� ���:�M2p9��[��3��;�W;�=Hc����a�F��B�C�c�>�)j6�V�2�U����v��p�Ҏ:t�n�,Z�Odִ�~��k[�͡�r����8D��S�W7���ѹ�QvѮ�2���<��A�#mc��(Hvt�U��|W��1�j�o`U͕jek�3�>w���x���'�$K��/�hm��z�)W���_�������/l�n������3L�2�t�����=l*�Q,���m����Q���F0A�����'�p.�޻���M��_����dZ���G횚�**v�@��SkZ�����-��!���`��	�\� ��x��|4�Q�j�|�u\�p���W^y���L`z_y�E�%��6������z#I���B����W�F�<61��zôZ�~.��>z����5����g������`g1�L�]�TҶQZz�j�F;DC�G��I�dk:���.`}m��!�d����?�=�#��H�Qo�� ���ֶ��:jވj��z�.�����@@W}���l��]��n&P���[�kݚ�n�P�q�vϥ?�����b��rѶ��xNɵu��,����6��Ĵ�X)��ܱX��%�$Ev�o���pnq��6�af�ǭ�$�G:��Ʀ��8<X��� ��^l3P	$�)����u�D���=���(\c$�Bm1�bqk*q|*"�����n���:�{7?������,��|�"F'Y:t:z=!��
��J#Zv]mm,/c��m|��r�}��9��MT	 ���*h����y�>��^�H�1����8uu���o��?��[x���q��s(�7�}��t��#��.G�'͙	�)æq�3��:����S �,5�H�CG�C�t���6��?e��o�gwܻ�Q����s�E;-��]�r�X�}��}.���p�ж|�����v�ɢ�.�H[��6ODl�xq�����0<4�l:g٠��);�ݍ����x�%SÜo���3Ѻו���Hq~f�3��e:wԨp�I��9q��8~�;����E�Ϟ@�k^ u�s�D@��|�2����7��Q"�_cp<v��u[��������q���\��Eᤨ����fp���Ek�`��h�`�A��@�JJ�
%�]x[|���1�gr�f1y���Q�1䱬b����8_�bT��܏h��X�r>o�<��?�[��"5=�sמC|l;E�o��ѵ=/s'��3/�"6?��O�d �u�Z�^T=��hB�3�`�x�A�`��8�p�ʍ�\[����{i���a��9��9ON�3�,� (�$ ���e�4M���]�%�/��]�˺�\�d�]*�!KE� K`��؜&��L�t���9'��|��ҋ��Dhz�����}��sD��ty��p�uMg��D��XJ}*�� �@��G�e`�XF	�!�C��[���dT�T�s(���ڔF��[�C���OsB0�8�/�Y�Y�^1;���=9�ut�Kԣh	ñ���.��މ1n<�Yb��SFL�����1��a`@S}�J;�ԛ��x|��g��0��l�̛�d0����Q�b��r��%�ۦE{��YF�s��fq�=|p�Z��0��7��^�Z�\��M9�#�6�"�1M�a�`U�m6;��e���@2y݁��č�����	G��o�^���1��ƿ�	�1��"!w�i���9E��,��������锩2Lg欧�^;D*NpP�G��.�tRw>@�s�W�x��?����{����
�*�N�L�CD�A�[�[���{[��}� �<�
����ᵎpw�`��/9�.���v��_����ύ��[�s����8AmĚ㕩:ɺȩ�!JD�����;��=)ʸ���f�x���݉�����8�_����D|2O8O�]O2:N��Q89�9�TFY]���d1j���QTZY􍻷���HW�����Av�O�C`YC�X�׿�tx3H��փ�l�����C�>��N�Y-`t�a�&���_ӛ82�fq�yaAM��@2�FBD�ۙ�%T6����%\�s�[{��%�������ai1i�������~|������;�{�Wlh�ŵ�JD�fq��%�Y|�gQ�n������?��n��&(pO(��O����������ҩ�xc\�\}�)#[���FR
��cue��mӳ�>к�W��d]?k}��QY�f��4��,��:�T��4��Μ=��)�s�^0�&޼����k���Ƣ)�`+S��( H�b��@�{�3le
UBӿ�仛��nݺ�ٙy�g��9iM+s(���]�֫gn��7;�$���k�#3]��B�������d��O�\A��H��XU�Q��ˋظ�F�}��z/_�q]Lq߷06Wb#������w>��X"?3{�ke�'.�ƀk��Ϟh�� &!�:q�����V�rd��1ڐ	�dQ\��y+g�^?E�7�db	�{��X�x��ȭ�,��������a�A�(���eC5�;���J���E������^�l#�S��1�#A{_"��_����e���1#�S�p����
������NL!w�b��u�Ч}��	G�"�_C"=>��e+'>]e�+���xF�{����I����e�,[���#(��̠����4ڲs*�+���O� �&}c�p�y��[5_$k���9�.׏t�x*���I�*�����#����k�ge��{h|���D��4�(�?%��]��J���|�����Q�s�q������S�Tb|��;uѥ����h�/#{�`d�6���ڝ*����y~n��\S4V��q#�>��A�aB�����[����5���!7�-�E���ݽ��6"7��l�@�oeD���T$a�kR���F�6@���d�ڊ�}x��?F<=�Hh����6���_�ƱzP���~3�i�L�OѲ�?���dFە't�j�VֲV-�:0$Y��1�"w�A��Od��M���������>��x�,�ø]@����ț�/����8��>|����x�/b�b��to\G�7�%����WVy�+������
���n޺n�M��f�kSj�`��a�#O�qD�O�I������'�~�u"��q���F �dX�NA��D���'�x��$���q����������u$8�#*�D�2�����om0����:_��轎�7��:n޼���XF��2�����th:俆�g�������sԊ�4�3{��p��ޙ𔾷K=�|�}9i�6*3�s���5�|��J0�A�A@��fn��U#�k㍷o���Xs�)�=��n�H�zh5��E��m��P�!�V?h	GC\��4^��O3� ��6���x����{�}��9�ǣ��M��p�����A��*r�m�sox�Tܭ*�(�����	o5��B������&�~/�g����?�%�ժ�K������<33mk�Z+�s�k$
���/�H������P��d�>�,vwM�dmy��E����S�N�ɹC�>p��=��v�i.��`�X60�,���K�����KW.)�*q)��?z��L:n���l����o-���>��V�e�D�3=��l>�oq=��w����Oa�Q[u�Fml��8��� � �J ����XÕK�x�{X8��F��B9���94��n<`��E���C ��6171}_�DL�;�kbjf�_�<"s+8w����Q��E�N,��Aig��m]gP��]�1�݂/<��[FȮ�m�8>w�6�j�𨿲�Z��bR������,���r���Q����q!:U'�<���4�]뻱[.�'Rl�J�g}�^���i�ԓ���z5�t��|��܏��� �ÀH���gl�$�Deb���[z+�<A�5��E�fH�n�� ��I2�L{'Dj D�p���mC'��ġC���-�j=~ʑ�2�á��c�-J"X�T`��5z�MѬ�q<��5ڛ�ٻ�q��&��7?����ী�z]��\��g��3�Ǡ����NIÐ���.zO����2���K�ࠌ��&._|�e,ͯ�u��8��G7p��;h�h���؆���(�w&t�Yd�H`1��cuz
�3���=�)T�إ��������B��ϴ%[���l��g�O���~ә(^�kK�Gc���D4��l���洯��hԍ��>b�ֵ��;�sq(�y��&��j�vwl
:��G�q�N���s׬���W�uX���!�����7p��5ӼL��ܓ���_�L�Q�	W�*��.=��]���).#BG�h��o�>�y7��<��Z����L���Sܻs��+1S |̿1�7��=��'�>-��@��r�Ĺ�O���݌�U���E�^���i+���ߔQ�g*���g�h$HZ���;�4�~N�9;��*3�L�m�/��y\y�2��y~|����5tp�2]��w�x����F��~�w3¿t�I>4vw臱0���+દN;]�2\?Ct��z�LMIg�v�8��|���Q�lT�s�>��s�Jx����DO'��^��~FDR�\_��l�厸��\��j3�h���2�>����{�+ʢ*A���#�*X=yz�ӳI��E����_���y��-ܹs��S!_溿OP�g�4�~,���,c��x�Ds��]\�z�Q7�����q��q��(��$��O�KϿ��g��j8ܔ����y�a��-�S�V.~�h��'c=���sF(-lMt�#O�'��'._��S�EY����F%Mb�K�f�����7n�p���\��o�e��K���w�Ë����Aw/0�����E�)֏���͕2��23U�u�a|~��Z�}����U#�Ƚ���<n~�g��٠����[<�b��w��}k��F���c~�*F'{�}��1�s�3#,�Ρ'�� r=��[a�B�nI1����]�Ʃ�\qڒX�+3�wЋF���q��r	��S�(�m��X�G�޴*���>VV���,���J��kk��}g�x���7(Y����je��v	�S��Y��D̏��n���q>q��m[CB�f�јS��aUc�b�A��{}����f�E8���f0`h+� ��謟�M�T1�i�X,�L���y�0ZL||�j*��v���!���wngfE=|�=ad��r�1�>��@��X{��IԻ%��Bk3�C���`�%Y������2%�$��H!h,���C�oA��Vh&��"4,<����||&Ph��|RO�t2F(:�	����Fv� �5�H৾���n�z�����?�G�,� �w�xgΜet]!X�!�_��S	�B~S��1է���yz��0��Qޞ��h����Ј���T&�f��(7l��xz	���shg����3?gN^��מw�~�[4�m��K�&贪4,t�K�T��j��؍@,�Z�@c8��1��<�����AħX>wS�y:UQ�0�o-���	�M����gPF�n���6PW���a7�H<�IWQ.lb�=�۷����h��M
Ń"҉#g��" &~�w�T���:����Y�Xi!I�z�<�>�&���-�v[�OwP*1���o�}#�6y��$�"V�Vߥh�77	�lzN��2����4��ň���l�s�����=��pe���$��:H"�,��yE��,]�[àѵ���� XY9G%e��n�x���w���V��ۿ�������'��w^��cm�ί�=x�mS<X�W��!"Ks�z&9�u9��׀��������Q"���L�\��n��^Bp�g��Ep�4�~K� AW�J��.\ŕ'^���9.+/q�����o����=�fq��3H�;�#�èe�Io���v+���]�U
�˲�1��2����p��<~�W.��g�}�Z	�R��6����9,�/�d�V�Q;m�X����)��u0�`�Z6eƨ�u��~�>`j5r�"����V�S���Rդ';�˴ʙ����
���ijAx��;��P����+s�N���ͻXYY%P  �/��w��3���P�k��Wv�(wxn����������	�
F�T$��GD9��y�ZC�#+��E��]���O�Q���y#�5X_]����%R����_�5�����.��wD��1��B*�7_���q��i$���#�ɵP����;�pY��K]a`��}�H�(�׎1�@a�!:��:�n���,��!mAI}�k��R��B������hӚ
���I���6��F~�.U;�����o���8���Lw8��gp���ߦ�la��������z��x��ό���w�/!�%��M"��k�ƃ�V����G��'��S\��fh����eZ��`�-0���r��}����d�$'��iO�e2���Ku�~�)K�ʘ��F?��#)��ʉub�Y?�x���Dy/��>#�f�f�`���@*[�91(�Gx4�k=�~c�	�"6�"�g�6�'��(�L�������v9YY�;È��V͖����vY�*�^����1�N���J'~eFs>>~��'P4qMLw��|����k�$WQ��d�Jv�Π�r�MG��k�����.�ϣ��t�HP�.�ͬ�,r�W�o�q
M���T��?�D�}LO/���	���-�	!�~O\|%iO���(#5�A4��Q1_8�͛D��>��8iQ�����(�����8�rO]X#-`e~e:�^zcF�9�j5��팬�����w]wƲm�H�m	�ťF�̯��Z+�����߳���5r�f��}��M��WD2=Bqo��%4��}\���6�q��*��~�F�!�FLOT�$9�v����/р���g�'(���������֓��{q���XlZ$��aXm*^�t7�̒2�{!5&���z���a�N�i�w	oE��ci<�me/���=RY��c"B:��ףfjE�ʼ�G=G�vT<|~�y��z��h}��6�K��JsR�_}�܁�7ʏU�h1���uwn<��_���-<|����W��(巭y����Du�1»|���xohY �BYB����$z�a�,�q�����r;���2��� l�� 3³W�Щ��r����-+�j&��!B�������9q��	�:x�g��@���?e@3R��}:�j�-޻��lomc>>�����u�~|r�&�O�^|�q?x��▒�ظw���|�pn/]�`�^�\"�5�J�G�����	����E4�r"���+e՗h:������|��Qӄy�k�W�0��*Y�B�v���e+-;--�]U;I��^dp�ϫ�p�S�C�qM���7����H�yz�"����A�׬��]�)��V����Y�ʗ�z�әY�gj�3�Zyd��)�;طIO?A��[66������Ax�r}���zj�_�ѷ�����^c�w��XB2�@<���=I�ob��������-��i�p`�&e�"u4���a��G�B��:Z���s��b�̀��z+�!��2�n�z������i�]!c�gm G��S�I�V��Ԥ�ʰk�΢�Ҥw��t��M������F�����̀s�W�p�hZ$,h�g`�l��J4�m�C~�6���bj�	y�`�lq��Ty�M�˔�H�'�;�Wo��:�>�(�\�z;���ġ�6�5���a��22:�?!�� �	����1t��ժ��v��H9|��sJ�C�Йb��>���x��i�p���ò�n����&�=���8��.�q��%0��e�ˑZ[�l�����nx�}�c������3��|LO�ge�b���k�]u�̺�!��b&�w������LM�u�������I0Jb*��F7��֝{��ؚ�53�����bg��d�D���x&c�@��Y� #��ŋ4M�[Y:�N_��h���a�:�t�.R��	=�[�ܩ[���Јqjf	�w?4r�Z��(�s�����M��Z������!#&h�|8�w��ǋ��?�'���:R�e��p��������Q?��GP�ᓍ�C�!�`\�#���yL�a��Hr�n�F��s��C6��~�{�F�������ls��yL����:>��=��p�x%7��ed�~�R4D�OY�Ti����:�N�X��m��O0&��Z3f�Z��� W*�7�m44�t�F�!2V�3�+�oe���jo7�(�����Z�#Չ6��ק@�B՜��o4B�Y����a�ƛt����w�Ĥ�N��!8�X����O���50���J0e01�T���?�a�"_��5V�T<H��������㎁B��xx��=�˅�Zh4���N̏�D�� ��>O� �{��Af��?�������}�t�WWfq��*Z=7a$���	Wc:��zt�s�`[�?2j�Z3��ه��ǆt\��	&c�6규�����70;����2��EloW��r}�hv��0���-bDg�2rK4�vq����[�w�@RJ*yL.�#�-���̬�)�e,��v�L�l��ҥK6��c:���R�q��9X���`Dp=�IK�q�K\���f���*A�����Νe@R�����6>|��$�[��:e�Uf<!W?��������8[\��nۀ�@�hh�YH�$�W��Z�'	�!R������e�U����~����;�_����F7�c���%���@,8D��-�^@��E�1�^�Y���[$�C�ԗ^������7�HPeVC��Z{��3�6��҆--��?�#�^��D�&�	1�����?�G,�B��Z�ܡ������r%���)`����1w��ۃ����J��DN����w	\g��y_�o������|R=�긆4x�'0T�MTU�n^���@aPG�6lz&�Vu�����}���;=$��Ix'>4jy$5��]��m�z�|�e�<�	�x��������4�m���N�3r��}�7���\F'�X��M�	�Ea�A�p�k�����<E?��"���˧���!-�~1���'�
��}��?�r4����L��Ou6Ml#���P��Čm2Y6XA���S�/��OX��~� �&#1�8[�����g�:4����Jk1�sx�{�X�ܫU��8���w�z׮��|f;� �&��c���hkk-J�ۀc����r��\�z�Z��6���x�D�����KCd�S�����#���,�9���h��2��iԆ�R0�}��Ѷj9WF�'�,9��m;�y��Y�+3�⹔���$�ltL�٭l�8�0��g�Dh\��;�PiO��u7?�g�h��2�R�!���q�"=�j�d�Z&0�cnf��6�4���Nh�i��4����� 6	j��=ST�>����g/�ŧ3��o������|��ϣҬ�n�
�Ӣ�Qt�N5����8�*G8�!!T!�"k�\)�����&D#QD�t��&���,A����U��v���q���*Z�)��Rיf�B��p��~��.�sT>������T:���֍�yܫLKe�C��tZEr	\�v��p
�_��j��)k�5�WA�w��Q`p���l}��sӳBG�a���x�i��#G٥?vtO���#jl�~���\�Q�L�tjO��Xr��4%��y��S�d�����Jy��,n�������G��\�b8�J���� �����
�*%�\�]A=O ��?���؇v�듟�-�M�;��������XX\A���h2��g�a?�oZ�:�Lz�Qi�>����İ��29�pF�	j�mYMH�A��l�Zet��m��!��I��B�
5�y�8�T�>>�Bܶ��o��ZRR��d���?P߯���ׁ����7���~@pwY�T0=;g��U>9a��cN����'�S(��2C*++�);w2 uH�6MPy�=����E@�L���a~Nl���yq��(���Д=c���5^�:N�.q���56x�4P�I�ғW1����o��i�hڷI-"f/vj�W1Y/�oGjz��<.>�2f@V%G�kW	>W0�O0����yt�{���|�G]��w��@3����6�Ҧ=P������ǻ��c�/���>zp��Z�b\���b.y>C݇��"|\j��b>9����v��&��I�^���hI��K�Ǐ�8=���2��"������f�~��Y����D1����drX�˪N>� �[J>]��Wc!���u���1�
D����C�i��7Q���vNv���F5fӅ7�76{qM�p�����S	��U��pd���c�Ə�i	��+�����ۧ���q������l$ʍ��"<���A;:XF��h��{ܨ��/���s�9�B�7���m�x�+�x��_�G�4��Ѷ��*"�.���t��L��cqj�b'pX��C�|���mp����C��,��}GVluu��|b�dr>Ǝ�I�`�J#�P�f��*��hl������G����QI�J���5B*�Ĺ,�dR|��2���mˠd���L͙�Sg�pz�8"�zkkÜ���qk��p_~�Ԫ���+p�j��b�£�}�nu!0&��/�JC��J<�c�Zf�
�[��ӯ���Y:Μ��Í}��p��d��4�' .y��_Ե�[ew$�W�Ō��C�!��z�J
�G>��P$����X�4x�U�h�z�0����l�����5sfy��8v��Zw����ј����2����W��2?�n�t���Е�\�I�|&x����Wqx��T<`���>�}����X^]Ar�ADm;�4�.MG�	>��/�Z3�1�,Ck#�W%��)Gm�إ$5���A��'���Ԡ�J�q����UE� O�����Ç��%���GJ�Wװ�[��N�ԁ�7�0=�����i�=�8�#�st�E�s+�8G�}��T��^_�߿ˀh����5Wt��?{�ϼ�5��(�|V>�E�1���K�0��4h�)K���0�G��*3��1�3#��3k�p��es�*� fp�C�ŏ9�y� H�>E�2���wv0;?c��	�it!O_~���N��猸8ŵ�`󁕙O�2�ޠ� ����Lj�X4MO�R	�
��<;�K%q���z<)/{���x��gmMj\�Q��k��V
�\]X"0)�PU�!�C?�ϋF5���D&����������[w��d��ӟ�3/�5�S���	�剝��FΣ��&�Z��KO=�w��!�[�2�?An�\�N/c�F�@oI�����S?��t���r}�{p�A�e�i�)x�f1.�������qX�|��'m�F�R�������5�mdP���1������V��*{�h�ϊt�P��6��3�an�U���޳ /J@�I���r��℀�@]�6��=��5(�,��&���"�o���xk���vz<���MJK�]���q�(�t��LR��u9��!�5pzs�� �� r�f��*��{̆�Ч�3<�i�/�.��pe�J�]��l[�*��h;9H�Pf��>���_"�1��\�TOL��	 ��F?�e�94�:����kb5z��� Ng�3������L������2�fmHS�n����j#)�QY�6(Ѡ?B�W�E�q����F�3j3���^��F�M�>��Ң:�z�+�#:7)X����o��4m땪f|��΀7H�E��d���$�h��`p��r��=��;��UӒ�ɓ#��i�3)�
M��@�t��M����̨߱E�SF\���:#y�o��n ����?�\\��XH'����:˨љ�,個�]|��\�|\���$��I4*-�Dk֝&�ӫi$�QLZ]i�z#i:�ИKBQ�z�ښ��4�����9^y�Y��K/���So�L��\�^9-po�(Y_�$���WU�	�����k|��H�ϋ^_������/��Hz���J+�n�i�ZV�5�cea���<���<A������&�:�d���l����-���zس2�a�Q��-BǮI�PP��y��!��G����{����c	�8�`H�צ�N�Pn�J���p�̓�N��lXI;�Y(�)��ʌe�d�G�c��6�c�26��ך3�9��I��S��L�Ι�A��*�h�*H���U��=��w�mh'M1��G 2���1@�'h8F�Kd��T�0V���̹5��x;�o��O]E����;o�?���+������Hq�s<�$�!t��Z�ϙ�kJ ��P'X�6v���̿�k����Ѡ�H�EF���h"����,0�l�J��;�$�0ʩ�5S��T��'u�ٞP!9��k���*
jm��6T��(�����K�C��u�n|� ���6�d�ѣ�H��jq1�u�Dmh�R�[6iuuݸ�$o��.*���/j��#��;��v�����>����k}h���&����3�tw�Hpf-���N=i�,���q�.
�s(s_�5��� �nm����]x�!�g�F�r��g�9ŕ��w�_�,����
����)~���.n}r}�Z�#���-�-=D&����W �}>�ٵ�ܺ�b�/mY �qT�����V����^`?ɘ��e��N�xp��G�r��^���oѦAo�a�V�n���f����d뷌~(EH\���Ra��Vî������Zo����2 �`��s�r-���P*:J<�s˴Ca���1�˹i�Ð��8#79ή8�\��@����q�k�#���<��<�^��l�1��O���;y����B���������}��<|\>9D�o��ǿ;��7~:%�:���9���>��9�.�	��wO?>~��3�¶K�P�� ��V�F�������-F��\�	�}�M:aFa��m��~:���(�������6#�ETJ2�	�7�srf�:�"1�����WJx�h�?��"	�]��g23F��b��Y���^�x
k�*��nbi�,?E�SXZ�Bg�hI��,	D(�Ut,��t��%�&`:BȥL� ��!����ht*���7d�cc(�RE�����\Q��fO�k�՛�7;�%�]#]�A����kO��zٛ������t�q����3zU[25��ߙ�X�i�<j"��1G��0��T���P�{��č��]$���J�[�d��%��&:Q��^+�j�#�
9
�duiI|Mx�D��~;5���~tw=h0ZO���9�-�-�7Q=�!���K �*�
��������K�O��r�f�h<}4�]�B���(�(^I:�ݮ�\J��ޗ��B�ѻ7�#h�^�pjmٲ?��V�g�&i�l��A<�����l��	#��9��7�{7�wym.�ψc�$��=�܄z��h�r{�A�р'�5e�0����'=��ɉy�ܝ>���\�W�"��R&Xr�/�=k� (����TV:E�T�L�8-�K`v&E �:j���	|R����$��g�Y_�4��S��a��֧g���cc�eJ@r���F��|�N�e|jj(Uk�����ͣX����~�pG��Gҥ����KJ������|wP7ڡB�A���zQ	��v�v-Ci�ׅy<�ڴ�J%E �������~�̞D���H�A������E��Jg�L�za�g|o#�C��0����M�
0�
y�=}�k�dS����&	�E�-�k�{@�iRɕ�ߧ���n�K�D4#�K�ة㠼�dЍ�O�H"~� �[�/�\{鯣���KVUhT��?�gx���s���/��7�����R�f��J��(���.�60���why3q/�}���G������:�{h��������4CX������L�n���"^���������+��#��0�@@`��j�	q_�-�Qa��t�[�\�M��~��,���q�"��~e�ם@��� [@��Wm"Q��x�{�]����Nָ_;h��^��d5��3��[���t'�'���y� �
?��M�=��=�����~k�h�ӊ.�����Uo��?�q��m���]�Q.�|v��� ;�7Gp��h�K�_��_�;B">eYd_�칝ig���H|�c&}����]�ٛ����3�v9�̰զ����{�����Xo���n�{�������g>~�����K.h*7O0եa��h4ڽ��؄|a�7����'����'	<�~h��S�4��M:و�\�N�N���}D���4��93#�y����; �j�*&��Z�_<���,�je�&�������y^��6���"4zb�o@�aͮ���סa������x��o[��t��!�Cۈj5m6l�B�o�4UY1D'4,�~i�`* l	O��Ԥ'��'���F���b1oI�$�S���j��&����h/�v�K���s���h5����T,a�'��TS�V �ܲ�-��	���A��-�z���?l����NG��c�x�ZĀ�/����qv$i��J �s���m��z=�a��K�^�l��aAt-tB��8��$A��������h�娲o쎶�ۢh��)��a�:��kгg�ILWp��)�yl����QiKKv�	zJ�	�78?�@!`���:���4��٫T	޻֘�c�������"�v���}<����z�&v�^F5��n@Ѱ���d�|� �)�[Q���K�8::�=�A&����y'	H�6(�y��h�v�a;�vWz��,+�Mg��
G;ȷ�X�*�TԦ2��]�3���E�_z�����Ĕ�%?Ͻ�ީP��wLR�<�}�e�TP�6_(1�Z���zQG.G�F%5Mg�B�G���g̉Vg*�!hK��I��M�'��y��݃}+%��*8P)R�׍㒴ޣ�M߯�I�A$��z���v)���"4�EM���#0�;�^|��c�6�
Z��tci��~D�x�Z�&�D�|���������Y�"k���Y�c����������-C�<����$�>�+9�Zb��i���K��"RKWl�:I������+W�8�ֽm|rc�60���0��A�߅ե5l����'�A!W�vay�"�\{�A@>��r�B[��O�ETKm^W�/��܅Ul>�?0p�n��{�������C��@�{s*��=ڄp��8D�S��>vW��ÑQ
��d�]n���M4 ����Q�P`0��z�*}A��g=�Id��A=�Z��p�o�ۓQ��9������3�������3m�d�p�Nz-�{��قLf�lS�S�r�E���ŀ.�Z�Р��XMir<pb�}C$�o��e��&��X<��S�y5�̯cX��ƃm�g�����۹���2���x=ǽ鴁bƘ8�|�{�7��xN� �Jf�Dٍ���R+A�n�:�E��;�ag:���c�B��r�)�����L�g��@x�i��H��7`��@�����4#�p�gz�O^��ݽ�X*���n�:7q��ҡ	��
Ux�n$#	l��E0���+Ө6[h�p�͉{�x�m�O`�K���'�ӫIC�����%���Ǥ�lO��`���:|7� �nF��Cx��wp��ke�3�$��w]�^���L3���"���d���Ȳ	>F��RkF�*��Y*6�d8�Y=҇���Y��S�a�t�ϩ^��r�j4���*�脒�8�y:�n�0���=1���wr.B��2Whb\����K���Յ�>Su��	���YVs��F��E������ſ84'���)��F��5�M���D� փ �Q���硶�6GBn3ޑ@�� �� ����&�a����ʽ�H��c�ړ�TU��5�����3����*D��>�e!��gc��i 9x&n������U�j�5!��ݫpr�J�!�"J�~��z�T>ԛ�iy�qW<qa��DC����C�yN���x��#�����U�\G�����p���mL�_DG: pl��z9o�m�kU���+��2���hR7���M���5�q�$�#(�|��H,à�ݞ8<���eC����,�Ax���#������@C��,��� c����%��]�Á�çR������(=MW��M� 6=̽g��D,�&F �>�����+�R��+�m�Dt(�.�͍70?�h�^e��Y!��m�AР�@�ZD
���@�w�u��8S�^�B˞�"�6B\���K�5�!�ƚ�����;�հ�:c����~;����{�~K�:��Uj+��3m|��3�0g�9���@��X��
ƴ!����'�6�]~Ҳ������7៾L�5�?��?��W^��Zf�$���S'���/?����Z�R��:�"$&���!�u�z���U?y�-����^@����j7��k����3��~�=|��_��/��x����]C��:x��Z}"J��1c�:���[�H������J�g�������2�q����+�I��{ض6���k��M��Oͮ�Q-���V�E<���Z��qm���Z6�či�@.I��v�,H�T�UmޱϦ�5L��������F/�JF	�F��^1ؔ���/�^V�_DТ�	���ǌ���?�u<�l���z	��.��S�xw���}���bI���3��� ��B=�j/�4<4ř�`hA�Qm1�Sk��|�.Ua�}�C;3� �8�� z�EՂ���؆�dˌ	���X�Ѕ�?����z�-|||��g
��%o�,I���Σ��(��z���)]�f�����7�� CeV�d��a�q���DR�SϤMǸXm0�[�2����hu	D	�a�����bV�R�M�1H� ~�f�m ��QT���buqU:�d�^}�U���7�4�����ţ��<�Wq��E|a⨡8	L$Ra:�=��pk(�4��������:�;�H0�$]���u��9j�̬\��~Śx^�3��q:�A���{{F�,�9lzQ��WFt��!B��DS��n�g_��%��F���X��v*�
�Arv	ٻw�א�7� �bt�b�+�2o d$�R�@0-iq|����w��Qk�1'�9^{䥳���	t�bqA�ς��[��Iǣ�o����"䕲�@N����G��y�t�UvlJR���P�kdz��4Y=y:� ��]�ح2U��������	����"��#j�����h��F�"��d��Y�-W?�<�t�q#��O\V��G<_���t΁p�k���qxd������#��>�3A{��5�7����&f��X���E��C�ܲ�C��4�h��5Ѣ0��,Z�oZ�j�Oܴ�`�g^|���ɝA�VF\�>��Q҈+�W7?�f��fS��
�_S,�8�����̜M/ihC�������O2�kbmyG��ik���S�8vF{�}����L�*ld���W�wO����`)�_����yS�!�О;{괩m�MbOz����n˲��vs�+�p��\�,X�����*;uz�`�e�D$:oS�����W����5�oD�R&�ѵ�*��{��G��au�l��� _�m4+��MI�.$�<:�!��_�t'Q~o�������}��o��v�3�#S���2���g��|.�^j7���a���C/ЎJ���]^d��Bi?�>NOz�n����ʯ�J��{+2��B��؅�G�Op�K�`>=o�nW����V�d����ALز���й��ⴷ�N�~���B������4��:�G�qIk�#,�-b>A���F)�0mF8�#(S0�\k-��hg3��N*Z���8Þ����Z�õ�g�����
4ԃ��z�}ǭ���R����zEׯ��wп�^K6&����y�\�X\W� ��m�M��K}���I�NC��/�gҏ�z�Azɴ�{~�3v����~:�r�I�Ʉ���-t���_�ǽ�C���K��F\nÀp�����m�Z�
�'	��������@�x�~�^9M ��o���l�ȥ��+��A�&�to��mk��Σ8��ã&a�Ot 9��z>�ٙ(�v�VLT��d�Fc,�	7�H0���m��o 57��!�p4s{�c��aHT=�jVd،�'An�ڗ^����F���/����ʛT����ـ���u�{�:��q N�IuzEx�*��L�R*-�hH&�qӡ/�-"�NY�i=}��!�7.�{
�Q ���ᗟ�[�p�����
��}d.�Ģ��qcޟ��k��P
��G������&�v��!T/M�&���:��-��=�..�d=Fr����x���x��\��䙜q��0���3�
��i�}(��gw����y�ӈjC�mᐕjR7t
SY��y������O��'2A\�Ҡ�ۆř4���k�4̦�2G��v��U	W��l���b�~˲��q"0�M5�rȵ�n��a]:�q�����O���ޜA���%b��\/[a�����:��b�.��)�[��2���� 1��Y�M��)>�~����HH�	^�l��J�2V��V��p�d�AB�4b˭��������������]�Dĉ����Cu�>�o����7���G��(ZV�^�#�<�u�o��φ���^7#��QO]�J�K�� K������}뛒��s�����}�
G�#�lc� P
*�z�sٯ����i�W��)x	q/m�ư29��PC<��9���q&�k}U����& \C̤�r��K[��7^�R���?�l�����^����e-s8��-F��T�,�gcXZ�%P�0��\�m�ŀ2`�W�(���l�d+U�S&)ν��}��w)��@[�Q���5[���"~�9�:A���k�v��%�3_�Y�S����x����7���):��!����^���`ma	+�V����=\>������m�̦��m~���ۈ�܋!��ܶ���P4��נƚ���@����>�S���Y�]��Y���X�qK+N	� I�[@JJ et��-�:���t�h^
�N2�r�
�[���k�xk���'�6�+��P(�@z��lU��ni�	���'.�+�s��&� ��{�H�n��F���N@�g`c
:R�; ��b�鐋O/Xf�������=�����d
ݮ��'v{��G`�4A;�.�j�Y��� NP,2h��K$È���JFt����^k�@a���G������zM4A�UMQ��7=NNȶ����J�O�C��*8c�G��|��\ڢz�oE�ǡ�v�ߥ�Sȏ��|�=��C�M��ń��(T��E��t6t�}7��F�:7��6��4Q�ַ��Zy��E?Ν��#웱N��iX��ǚBY�D�Wժ��	h����ݖ��$`>�1���1(i5:�a���Ĵ�ƍ T��yI��i8�f����+�Q�հ����R�ʍ1*���u����<f�U�l���JD&#�`T<3�HCK'(��	�{�p���	j���׾�g�����I�$\ʻ2�[���>CpU�kt2z-�4�UYd`�.�,A:e7�%d�h$�ӊ8U`�=�5�n7�|&c�8qn���O�ծc�&/�8�s�G�&g���`g���1R��s<��>�E$�4~C˪�	l437!�yn��{WZ�������� 4�ww8f=JaF�ɰ�H�ۍ<>��6~�d&���i�9{�L�N�ס���T�h�������[Ut�Y<ܸ�5�Bjng����}E	9�@�9����H��,n�U���������VSt*�:�#���
�~��|�_�2>:MG
��\o5��~-�ܒ5�KM�	rྎ�~�}���X�Q�ke_|˙'�>+YU��M���s)չpi�*Ͻ�������6����/���u���i��^S�J~���a/[@~7�����=ә��t��Cː6]�s%A��3ss���/�������_���
N�9��=���#+��臯����3g������|��������#�x�駹���?��>��)�l<|�g�}�+�,0�T��Sx��,(�T���Ϳ�3�����޵��'��/}	����!nݺ������^����3��~�+X\>���z�?|���N��[Z��\3��Ф�n���@��_|�{/� 2�"��G[���U���܁n�ᩫ�q��7h�D>?��L�m���m�<�&� �VGGX�Y�Yݯ^a �`�o�����?��T�g*8�����iSY��+Ƈ���֣M��Tf�M�=�S���mJ�X���gL"��5�m�~���\���O�:1+Dh'j����zv=���yiWl��i�H��^~��5YL�zNL�^%]������~��?�{�JXX}�|���?����#F���L�ӨԎ�YJ�}���>ˈ{Ǵ�cQ-D��gm=���%Rpyv�`��D_�9|�^
���Q�H����8�"�$^�9�A���S�r��3��I�)����2�c�+K�3�D��k�j]�r+F�A�0����b�J�l�D�a�r�G9k��h*����{�[�գt�H��!����d'.��ZAA��A�`_����4�撤��@{WM�n|J�=6����1y����y�؉o|�g�(,����U4L�@�Sj�hV��u�f��b�Skum��G`ө�m���ڕL��X_�o�Uv����{t�Cl77��-�X��f��j��4�2����ӂ��"Lc�wL��H� �\�#�G%�b�ס����0ϸ�����>�_�e�JOpl��g�_F&5���׍Me��.����\< ��[̨����O�����q�v��^³_�9��7�h�����$#�o��Ztt:���&"A���Z�!�l�`��w��RE¬M���DYW����P��V��=��)������]��E��7�Ā��ղx�u��7qD�/������j"�&��d�=GH^m.�@��֨>@�4��<��I����2松C���Y�M�%������Կ�2œE���t�*Vv�D�=C�Q�����,�\������q�?�^~�l1�X� ���Mr���=o���3�+�t���u�1��z��Y�s�o�&0�^E�C S����TO4eε���nZ����X�C��g['H����q�~��(�db%����;���x����a�t fj!���k�$�Е���8�@f�	"�E�&��w����B%N� �!Ȋs�s^>o��n�N������yD	�qT���503��{�����_��X]�1`��[o�&5�E���O������(��|:�\�M`�f�ϭ����'�C��7u<��	&�&:�"��=Lztr�C��o�߾�o����/����7>�Zч���_����{7�;ش�����;���	�2/������@n�N������ο���������{Rd�3������� ��s����ğ���cia��o��/����L:Q����c���~w�����wP�n��4��:���i��IA����n =�B�������4\��,���YMm���ac�G8uv��������7~�ૃ�|���J��ae����d���ϠF [���ϥ�P��?k���~�2 va6���gl�#ε�R��W��"�A����@˭ʎ/��]j��V0�����w`Wp����e�a�+m+W��"8��cqf�o~��������*�����g�q	�V��_�&���h�H����=}5�a0��t�n����m\|�2�<�%�,�G;�AJ����D��.�KqJz�G�C���`��J&R��T_�j%�N�}��+FL�̣��~�h�ziX���X��c�=�,=�����C��i�{bO� 3 0�$@�����H˒���Z�dծe�\*���]k��j�DK��]��H�"	$@dbr��o�9�s���7�w.
5=wn����{�s���U�	GN8�i�rp��Lr}@����U�s�Q4���O.�t}�meih
�P��}�BMu��*Ξ<�Мu�
B���F��}���'�Wz:0b���B?�/״�8U��D!������%KL�]m�}P(J�V��Q����=�(4����h�����`l��ӓ~?C�Ǥ�}}�f�{ς����-�Ϋ��.���߅�ǂjm�:���RG{*�JjD�r��H�Nl�XZ�S�)2�����u`I*ߣ`e��MJc-(�?�bˮ�(�_���i~����?F��̨ݪ�At\]��1��f�H0���ݦ�5�:m�t�p��Ex=a���;�z��(c�	F��n�"��S�,�'$<�٭��	�p��<<��-tiXZ4J�:��`r�:�͎ؤפ�R��>��4#�6������0/d�£��M��D�R��=���V�E3�-���F'Uj������(T3�,�itl�Y�r�u8B�e O���65����  ���	Q�����F��E8�:S:����8�
�@X�n����{)Ӷ~~V�ۖ�5<�]}:&�˂SOL�̅g��(S�B������󩑖��a� �������n�dO��⥧��y�?��
�Q����T}�`�������)�� �t�M������iq�c{s��:������b�@{,x'F�a}�.2�M�f���P&(��]����0�����w1(N iAr�!A!��t@�I��<r�4���;)8�&Bad|��eb��:���;H'��ةsp؃�f�P�M�	��$K���3��\<#~��<}�,�x�E%�S�i�+��0`������N ���O|�5�K�p|a�AR�Զ���M�(;+�q������N,�N�ֵ -q�&���S���A�$&F������H����\�N��{����*')����٫��8�"�F` v���E�
��#�m�w�2:�Bf㉣8qx� 6I ���}��o�&ʵ.��?P*#�ӎ�|�5���c�)�ij0�� t�V��8���O}�Y�v�J�Cf�[���zT�5�E���_ B�^V�O'��ŌLL�� a��C��!����2��j)5� x,uZ�o��q>[B���k��Ε�����rF#*�_d��j�
H����=�\>���#���/1?T�M�ruć����ao���k/�wR8:��o�������OQ�1��آ=1 ���w�'w���}kN�&^�@(������1��T
厉�X�./�gH؜u��4�)[���Z]�6d�WN���Y3Ǵ>J�.�u�
@4�]��%�(ܣ(��U��ɅӰ���4� �b�|.�Qi��������x���'�P����^E�NN�Ħ�j�v�' ���S:�bb�b6�㴱�� e��h �6 i��}�z�{��!�"<�~�o%�~����%K:�M?z|���.T��-ǯ���<�<�e�d���~Ou:�����hH�K_I�T���yPy�����*#�*������KC�=��@��:�X�0:Y�D|��/LØA�-��}mnN��B[O @C!�N�tl-i�5��H�@�(d���b�#����^�����N3�����P܁[�B�Y`��-����.���QF�A�͛���[p�T�������k�mU����W���CQld6��1���/��;���c��oӨ�"NC�W�ګ��ޢ6l��WA�Ї�c��j�n�C������Rk�Ny����1�6���x�ZZB��+�ǭ�'�]F�6A�V�2���53)����7
 2]�����o���[��%M���bd˄_c��F�v��=�]��~B� �O�h���ib�=:�æ�RJ!MF��R2�n�u��Vp#�1(��
���B��H �HWIi-62��ԴAv+
�o�^'O���$��t�$%��o��^{�5�O����	�j�̶ݏK��32�n�}�� ����{�JCj�	/�*:�~s�/��۷k�ܧa�l+'Z>[a�eCbt�u���!6v�u��MH�,Ho���Ɲ����g||
s�O��袴��=��Sg?�{60�F�b�v���T��3gphf��G��$8z@�fFzwS	�>�fѧC�0wcwcs��K8�ϐ����ױ|����X?��_T[p��uDn�\���|�������5�356�7Do�?����[���&GPY%psX{��C�Z@��V�z�Z���2:|a3|Љ{���"նxl��*J+�#c�������w$�ſ������_��?A�C�]ibl8�0�t�G�u3�b���Ǌ���`��㼶=��w� ׃���`�f�s�p��"A����fiрM�X�m�T�u:�$0I�&pqw�:��<:ǰEe/��*���Ӏ��,��A�=��.�� 靔�I6�G�d���K�� ��ڿ621�ݝM-�vi����b���v�$h�- A�.�R��	ہ,�Sh�:�_It�ׄ��@mcym�q�Kz>F�c�4p;<��-�瓘��������^��|V<��c�Wz�AJe�/�9��O4�mn/���#&�(�`;K;�}q����w�������bPk��7s�,J��S��ZD~h`7H�;S���J>N�$�_���1�w�&�.�1���`\�w�^~�rO0�0m ����@�V*�!���n��uתI�j	�9������,��i��~�T����k�42 ��~J�}�B�#C7� ����=��Z5�7�QMx���4��~��Z��{�G��G��x������ ��V��hL��N3�ȝ���:zM��C#	�����g�-�6f9p:t���J�+�!�^:�#%=�с�N�ַ`xX�|�t-D����8$�l��\.0����t �To<1����K���9�d�M"�YF���5���+��^�2�ABU�M��x��Gq����m��#4s�X؋�y^GP�v�4.�pH)5��{*\/F����l���g�!�$����x+�R嗱�(.^x�t��S�5:�EEå=*�0��EM�aҗ���i}!z��ib!���T�hi`6JRZi�Mx	�-��-|�.�概;��x�!�7+�L~+سJ�����4ؿ �6���c��d��3)Q�LӰ�����aQ����������C&*lIEԄC�K�K6�ͽ"߿T�� b4��t"��j�8�\Zx�o�^�hv4����7����C:&�B�F8�?���s?|���O}
<�?z7��t"6��*`���nP�?������(��>X��R 
DPm705;��ʛ��8|H��
���:%�n�ck����1���>������UԫE�'?�g0ܤ�/�4�UmxM��ɏ�{u�-��L��&�����<A��/��?��_�;��������%:6��s�����]up�萂B��QCf��u�vj�u�u��i<v�0�=��|�/4����m �d��RÍ˯j (�"�n�I� �k��>R�:@�uծln������ŵ�V+���	Tk��M|����#���hЪ�Ź�~��wP�$��^(D�$�ớw�ڋe��g�Ye��=�C+�w���/019�"m�d0��	JSX���C�6�����iՁ�Sg.ⱋOs�U�֏��`w�Cn^k^KH�b<^�+��3�3�����E���w�Hnn�ް�@B�ⴛ���Dp(�ը��1��.�k�^�� Gd*����B���R����aE��Xh[G'�Y/������(��`�lNi�Z�|"B�����NO��v_���=�MG�Ťz7�|&�C�Cd2���ܺ���ON��m���D�WJ���2*[4j<�|�b��Z5��>M�{ǣ*7�h�i�*��;|
����e�
�I2=/=�2�'��OL����j����(�J��I༂T*���q�K9%��lw�v�</f��`��k�r/���!ui���H;Z]��jʴ���Ra�p+�I3��vc�'-1�5`6헓�chD�����(�rQ)m�}�e[�p�.;T�A�vtZYI�a�佊G�G���x=����fw�{��2����NUM�K�R6���ui�Fv�������T>�~C:K(��ՑfZ�^:�&O�iW&���@/=A�pv[=�	���H'�F"��ډ|Id��� ZiHz݊���"���t8�	`rd�_��\�&Ν���ͧ����5���%0���^�g����'���S���T��\j1�����Q4~��VP�8v�(r4p�
��VV0z������ۘT�K�x�8�z�M�s�.��B�����-�cA92���>K�<�}��i+!�� ��6������e��4�[W�_��אD(Ռ��H[�fo_�݈�%�&Z�֖%�d�+�i�����ݧT�̢ٚ�����3�T�|`�g�}q�6~�$���t��{�3�}nB�]%T�ώ�x$��A�}�ay�`r]cj��gh�H#w�F�AC/���ġ����8,�ݐ��M����t�T1E��-vC��2bȬiY ң����&�����v��.d���6V	��X8r�x�142�_|W�����{��i�M��;u��}�d�>��a~������X������w0QC4�X��C�.׹�B:�OV�8z�u�¢pS�I`tf
�d�A��P �8_�q����3�oҎЉ����+��T7F#�k�}��o�����jU��t��~�L�޺y	~/A�64㥯�g�z���b���.�Y��ԦR��F83��zxq����.a�s.2rf:���1d+y��+@y��4b�Q�L���h��\��:��ݶv��@�-̣�]�N�!�KE��y��U�-Txμ���*���7��w�i�/)��ݺ�^a_��*��~��:�@Ď����NY�z'�R.�%��T�����]icd�b(�RŢɉ)lG���/���+��[Y�¬p`�b�F����N
�,¡���6h��	���w\ˠ�7���l�.#U�f�Ž�.a,<����JN3c�s��$�2)	��f�؇"�]���x"�=_�,��H�j�fl�'��=v�jW���~|�q��2�Q��;�n��ݵ=^g�BCQ���w1�X��{魇�;{��.���U�T'��5���F���x�o^ն�&�Y�DIHXj�k)��g�J�`�2��d�)A`]�������Cl w����l������niP,�W��P՘����y�Ǽ��Ņ�'c`��H�z��A���>(��K����~��}�BG�a�% ��oh��a����sP����?����T����j��&�:�_l�K�%�[���uzj�|�l�3�\!�R�![z�E�k�v�����	�.�p�^;x���ݣ���/PX�=��$������#0��Zhӑ�,�������hJ�PJ�|�C��Ŭ���466J0VW���yU)���r�,���;�Z��Ӊt�� ���k��R/��j![��!�)7k��!�.�'����S��x<���(Ν}��~��v�`�q�r%C����D�������b���0���g"���Sg�:�׮�xa��y���5���5C�����ii�o�~#X���\:���TZ���˸x�"~�g����t@*��([9���Θ�����&})�J���,����4�5j� `2+���ZE&�Xꆮ�p��쪾�����lJ�mV�f��h@%M�Ҽ���`Q�s�������*=���,�`�F[~�� 'g�49xȵ+�2O��M)���4�2P#��z@��_��*���Z�ݜͻ�q�M�fT�\�����w�k�g�Zڑ��\���������pt����_��_�pĳ�>�/}���=����_����&�_ss�(�*1'S����}��lll���L�l}�3��f�FC��bq��3�5Xn]���I�e���K���)�=,�?��Y��E&�V
�c�F��F��H�k�zr��raA�H����g��A���de�����Ҍ|LMĔM`��@v�^x��f�/��D��Xi 6�E�o���CJK�����dv:����X<2;��a'	��=XB8�=M�25��O|�SHf�����hh>tq�r3���
<����1}z�n._�1*�*��&xicv6��'���}�;k���a��V���j�z������l<,���
{��1��a,ݾ��a�lK�Gz�l�1��v�J�~	������I���)d�s�:�	k:�[^����s��w�����q?�h_�T	g��d�M���>�gl��zV��b}gn~g!��L�)�!r�Q(m�i�d�a���&R�M��M��I6'b�m��yq��F�0��&hl���r����r���U�hV���[F���U=z��.�9��φ��m4mi8CS���f�b	���eJ����V1wV��,#�V�	$�%�A��J[$=s�����<�+<[����xծ�aS�8�ڔ��;p*h�g��t�6ާ0,���r�ݼ���,�|A�O�]�^�uҦ[��v�7A�T'���؈o�	�7��Tĸ�̢�RG�) ���lj�C@�L�+�~n˾6�TGdpƢD�±)�Q�N�~G'�%Y�o�0��6-�5���D��V����@Q���4$&	�;�\��?�+|�xߏ�]>�u�B�e����Y(�v��tZT�A zt*�n_�=%	#�T�A���rd(d+p�<|���h2�+�]"�尋WQ�Ճ��p��a[� ��t�|Ie��_����m1z�I��N�R9;���:���F�ȈO�Ƅ&��)Иw���N�g>�iwpj�r%;��F��b�j�ӎ��Qܸw{�=�G���yV�c�Bhl�j�ҿ�tc\8�B��@2�&0X��O?��o~� ��
\��D�=�b������O�]L�Db��4�K�H�F���,
���H/��m-�������oL!/��F�Ҵ�;0@�`�^����&���HU$���A�,�����j���3����N�A�_�2�_J]M�!�d�����zm�<'��6�.I��"������[�'ZW����,��?�W�:��`%K�uRT�G~O��V��/\�b����'�������w�u�����_���o�~�g�g��o��J����!�Kc�5���!�g�Z����OM����r[`v
<�&�Q: �'�l���:���0m���2��H���mX�ocȬ�X)-�=����Q,��Ux���FD�����7q�����[Qi�m!�#���ިz�
+�u"A�N(�����3�RʎdV��t�U��	T����b���\#�w�n�fP�%���$���)Ϥ����%�����^|$��wn^Ghȋvq��!l� g]�ܬ�|A��X��ô����&f&ao;�Y!j��P��q����q�[���p,��/]��h�T�������FƂ:\(�-$0=��Yݰp�T�^��c(F�=ܿ�f�F".�{E�c(�Δ�YOO��"ը��L�?g$�xl}a'���S܂��@q7�W7o��p*�x9����%@�lM=��d�x&qJ���4�rE,�8�Xȅ��[\c3FC�9�);S���#��	x�8�ۑ��5�ܟ�Ә�� �F+��W���ǰ�I#����@8���;؏!���+?-�c���f�3�W>�?��3���ǎ#�� �kWPK�����r�+q���t�b����m�ie_ }��������M��si����	�x_�����kq�9���=�i���A^N�w٫B3��-�5�'�	�X[�ν�G�[5$�z6AM|t��ڼo��L�dpF�x��}�Mi����<0�E�FJ�fF�vh'�ʨ -�K���r�(�����O��+B�w+{@��)�5n{�c�J_7�2oj��ޯ�Xq`����A���qK�$�����F�G6��k�ǥ!�V-+�4����$�
���h�+�9X��>����G�S�V����0�n�E�����*�����l�azx�����#^��� ����!Xm���������̨1re7��:��8�x
�����g���tb�f `06=�#J���[�aw��������8�gC!$�UɤF�Xm��Fݹ{�����/~�����m�����IS�E@��x%��hY�j�铉�F��O�]��%2m����������̦f-��� 2���w�G����S�"`I�M��S��6�~OS�}�7PK���M^g����������¾F�<'�"��ej��#�jY=y��/ҭ�0�b��;��P��F�д��r��#(��Q��@~M�U�_�\zm5���lRצ�	�є�O)Aٛ"o��u�P2�^Dy�'�
A���!�NMk?�������O��\}©�k��k:�<??���=zT�֥�a �pST3>��H��㴽�=#�fw����ׂ�gDiz�:D#�<�@�5n�$K�� d����М6;Ь'��������!�u7�E���N2O�9>1�J��!��F���z�I�|+^]�N?���U�=a�k��m�$��l�E3)v�1!���ԉpA�J'JpЋ@ԯ��ҡ����#He�L%��;1=D����v#�*�79>����!�L�6#(en��^t�D,� �c��ˈ��<�m��a�t���yl|-e�I�1��vS��+e�:u��v����A�G�I��� v�7	y��F�Qf�13�V��{l�i�Y/ot>�`wl:� 1E`���i�D��&J�;6y�`����	�G�x�{�#N�u��ǽ(b�\��;�\K����Uxx?���^T�T	�Hd�Ak	w�����Đ��m|�Rƀ[�iO.�#/�4��x+�Қz�̮3�b��6Aj��v�܋�.moW��6A$���J)ԋHlT'��'��}�*j�,��-:t�/SZ��	7��k�QZ����=DJ\ρKt�mZ�e�d�v�}p(=�B�R*�l�����a�*ϼ�a��2�s14�{gB��R�Ma�`��àɌ�(�d����C�#I>~p��.z��H�>H�K
���5��K�ea���L�o(�E��ﵧ��I¬�7��$��g%��r�Jԉ�șE��.���pJ�[ȷE[[�K.��W���j�@]*>]���J�00H[N�����.e�G�G��x_��#h�o�2[K�eHa`�);����򈜗�Y��GG&U6�I��!�>�ɉi��I^��o��0�p���.�nTh�Gc1:��	n^���Y>�U�g�!<*qe����(��z�P)���A*�Erw�N�' :�՚*�gt�@J`�(#A ��,�M�H��郻w��n4(��"p������P�4*M)��4�%T����j�F�mfNҡ�E{�|GK(�����^xAy����J�;M�v�����Ry��ߓu���Ū���L��@�����HYF�xdѤ_O2�2`"Ϸ	��ł��I��!���ε>Ȭ)+�͢�`yH4i�t��l�X�3�}5��Ag��܎��B������d�HV��������Z���OB��#�'D��C�Y"���k�g���t���FfS�e�>G�� �(? X��jp}��*����+ͅӮُ�(ƈ��]&������ą�;��ӓ�����~���/������_����/�U|��_F8'�K������X<uZ���:tt�RGN��[bT�v��	.��൹E=Eh��9��^�N�@~�G��Y9	^{�S��k��E�E��X�{4�v�l�x��'��#� Y���5Nt��^�@h5�^��)�����!��cbjk��t�~��1�S3���ۢ�F#�k��T͂��h�Gxo�J����u��1ac/�8�-8�b��0���Ȕ�SE"��`���[X8M��o( s��IxFX�M��֍�*�'�.�L��g�	�"޿�%���G-x�)�u��ܦ��n�>n�~�k,J5U�,�� �V���,_k��g?�7���w�b7�G� 304C{dQ�>�ý�SEoąj������]u����&0^��>���k������u|���`smG懰����^�C�@���g�*/i�`wbt{��V_FBA�	�G�Q�exf�p _8w���5O�#>�9[f��J�,�0&g�v���l�ڡ�f@���Ti����5�16w���{5U�����S(�=R���Th�켎��n�x'Ν��}�ȧ��Aw���p����TXg�x���-�6�$��B�-=�]���[!����Q�l9o(�&��jQ�a��'h�>�*��<:���]�m��Ā��т���ajq-��Q�J\G�G���F5Z=g2��h��+:�}�v�k���ދ�7�E�Ρm!�W-R��a�rI߰Q�=)O�mn��jut��Rw�0
9��ښ���l� �ڣ/�xuM�����֩�Ar�i}�{���A�;SHp��pX����]l،!\F�b�S�ٗ2F*ͨ�E2M�6>���;�i���A�&���8����0��*{ת7�)
o�@'''��)�t�pvl�P }:�X(�4�����G�Ѷ$p��W*ӡ/#�ڛ5�:9��/��]{��/-@Ui�5�@�@CJ ����n]e֮_��o�a����Qt:�q�:�F�� ���gN�L�^���jx������5|�������c�H&�F�U��$
��*{�L�f��ڇ��A���,���x�?����7~�9�R6���u��=�+ _�~iY�彾�f+�(��^�W�FLV��@R�idoH�]lxX�p��k5JV�(��:�}6�_
�\��0�ls(@r])yko���I�f(�k5i��I_#�u�7#�v�@���uRO%�a�g��W�E�m��m���R�� ���/+=�B�}rq5�kW�(Ȝ��EthDK�����[|�[�Ɵ����ǟ������?����Np��>yJ��e�E2�=�@����s:�	)�=!:��I��3Y?{$����KH�n<g���pC6U^O��k���J�M2� L�1���O�y���$�b�o8���
��&�����r��Dq��K�q����p0H��Y���NU,��*
\��eX:YL;$͡�e�8l��ß��ë�S�{������Y̞N!<<�<}��o`vbN�;�w�ű�&0���ar�(~���t!<,.:IiO�OH?+�<�'/|9���/N���94�;���!E����1���?%io����X�5�������j\�z߉'�=	�K4���W���ϣ�� �����x"���?|�[��]E�ʀ��;�s�m��;�ʕ��t�/�F�V@02.�tp΅PK�v�*���Q$f��l ���E�B��5��v������HVz�^6�c�	��7"(`ԐJ�"ÙSga�Ms��p�F����^ۺw	��*��{����%4m�O:�384S�́T��i<��Ϣoa�R�¡#'�[y��=��37��B�[�������K� ��843O悷�♧��C��F���J*�o1޳=.��nݰ'�~W�Ħ�$	���'���F�I?` ���{������xߚ�&��F���ŭlR�D�J�ik��c�72�� Ӭ�rV��>��L97E��d�	���@	���k8���f"����}�+b�E-�Y�QŐV-J���Rgv��R)i����Z�����>�}ի�@���z���~�G��xߠ8�Eڟz3ќ ��)�N���a��L�*�AKϩ���\vQ����y-��g,}�Pc��(2�uɤ���&�i�j��a����,|6#/����������uB���9�/�P���!:ь4n��:��k�akw������JZ
�{���,�^�޼���Ȑ��T�R��`Z��L�$	`Oak{VWq��c��r])yon,#����Ԯ*����1��ГZ�-f�*'­�kZ2�L`[ub��K$J,�� ��$��I���Q�ݾ���U�7\��Ųj���@� S�}���H� �6)�A]c(0�~VΘ6z�efXK���T�*C*��`�l_����m$��]��Q�x�����
}�K童L�0�YuY��DI@���(��(X��m�'97}����/ QJ:4��f_�r���&>��	�
��9��!ɢB�A��	�@�9|X�%(�~�2FG���N���ş�^��p����=�Q�	0������h��f�\}jr�R0Etxz��8m.����Q�#�1������C���s��pHz��F���Cl3`@Q4�!mlOrh -�[�u�I��]�S���G�����A���i��#���� u�~�fƬ(o_F.]C���s��K��ژ��_u��[0k��Aa5'�o5��C	�I�8�Lf(Ux��Q6y�CA�Ւ(�p�ɏ#�� �4���C������Mܻ�.���>�gp��GX��In!�`o�k'��\K��,cG�(�[5����L�2���w����+H�y�	�<�%TF&9~�����Ƴ�Et�<��)o% J!4�uX$�ꖴEF2�a�������7�
MkS�#�9��V�x�qï��=\��Od�`=�>��[����Y<�۷���Sgd���0�0�g� �y��;�;6J�8<$�uC-*�|�љ1�G�ˬ�,���={�H-�@�n�'�K<���^�/b|({�$V�]�����Ɲr&GA1/�tՌHp	�ӡɣ��"���b�=�X���sŽw����
�<v��ı㓪y<3>�nN��^� ?��/~���H�+�K6Nd/�F9T�KmFi� y-#���,�+R~��&t@cG��gdS�t�:�����=��t���7`�R� �0�C�k�h7�_z�xd	.+y�
�����Zuh΄��
�N�0�즖̥���32�e1�#b?��[I����O�hW�Ny��t��v��-6��w{�*�$��ʲ�#v
`mT�^K{� ����&��q��[S�Eu(�(|�S����<��Y�Mm�?y�uj6�v+�}[<�р:N����WrE ��"���qح���d��A``
���(�`��!����+أ����xFc!�w��q��15*�<��.]��Y7;��Q$�#�������}�[L�O`e#��%�"�k��$氼��W_��_� ��A�G�9�h����!�"�� �(J@)\r�$l׌&e:�Z���1o�~����_��_�'��r��;��t��o��t8%�&���
��ϼ��'�[��=��g����6�H�S�RB�����c��#�2~��Tt��Tl1�bs���Q�ie�5��g��If����g�j�*��e[�u_H���~I\�A�d����x\�-bL��]2�WR�ղ���ܑ����l�_�d>K�T�bL����+�ף6��%�����=�M�!=��^�0п�5	8ޗ^zǏU�>::�K���/����s?����S�,X�O��L��2��?���a�����dع���<Ət:\����sd��~O�ʎ�K�e�ax��ӡN� e�Q�rS�53��D���|�k�bou��+��ͱ�!��5��h��6���/����mT������{�j,����c�u�:�^��z%O'���Ϗ���^��vO�όs����-�/���n(�r��Əo~E!��=���SG����N�jy�Sh�
��p⢛;ą6��7���X��".3>v�Y�x�77���OK��:�t5s��{�Ƈ��g?��Q��Bu	NO�`?�O�ܮ*���4�5�E��:�~��ӊ��jD[�ne�;O�j�s�R%�����Yv*]头��h�i�[���`��𲵁3GP�}���1�r�����%�"QfN/>�H<����a�'2w��E����կ}�k�4�^Ν>�W^��L�L���IL�Π����^������H�1��$�C�>w�i�D�@�]�9�i�~,1N ��;B ���5j�:�w�N���{�oQ�gK��|�i���E=�gF�� ��6mp�h��ť��J�$Z�<�m�(=םFӠԒ=k7�\�&�����m�-�{��Y͢Zn!�g�|�J��A��d^��az�Ţ^�+Q��j#xg� ��|�qJ_��g�"�6�O�0��"�P���a�߮@ȗ���djpiҶ��?�>0�(��I{��ե�?����Z�
JF0B��� ��!� �=R�͑r���T_#lZ2����h��L1������ǣ�y�O�;���ߤeB它��`)2!�Ѣ��A�;C��b46C�P*���#*u����"#�χ�P�4=���&�k<�2}ZC���tr��4��0k��HP5��c61�͹�v���ئs����)�YZC�uj��j�~�}���o��<�~�_���u@I��n3
�{x��?����h����i_O�Q.�z��S��Μ"�c�aw�g	H�a�����L��i���[[���|/<�\��c�Y<�H��۷nbiiI�����h��0#��򐲤�.d�\��V]�D�ҳb�#�Tj�hI�Ez򤉺\6��4R%���C�ՠ�9 _^��F�eE�V�(�^�`�g�f	ޔ�=ж�qP����]��D�қ(�R��\����	p�R�������� �k�L$�s��A�-���6�:L*�Z���I�Z�戟q0},�[�.k+���y��u�Q^?O蟱H�(���w��Q��I��L�w��qs����Z^���b�1�����7��?�<>��G���}C�.����:Ο?���
ކ��l�E �V�E�{LJ'�{L�^�[Λ�=^C���Ƿ����B���k�}�F���ѱ	�x�P���C��'�%6�UP�՗���~�#�2Y|�?ɧ��~�u����R�}�e��H�sX��@#޺r�|��\q����
*�F�	�	P�>y�{���{����7p��e|�'?�{��lf<2�|>�=VE!]Fbz[�ظ�D�� O?�1<u�	�'����U[�L�a(� � ���ck�.陵���T>���X�<�x~���t�=��994�k׮)�8�xJ	�oܾ�b)��s�u��5y_�ʹ:c ;?A�N��Aצ����w���$ #��cgu�����1~?��g��,|�>?��i�j���Z˄��	����>������{x��H0p��D��(��%���bbf#	&�N��_E-E�P�ũ��X�@�ײ�׷����~]z�Uޏ(O�)W)�W�i�p��H�FƇf��k��~1��F����/A����kF�i��`�� �թ즰�w����|c	�Hm��7��f��a�8v���㉳�^�N��\!�4���wp8Wç>��*�ZnT��Z�}p�ʯ������IO�U{�ѳT'$;�c�~��d�g`}��FǦ��~�����c�Y��$$�$�^�'��	�T��K��d ��S�=;y���kNsW�V�\L{�Y>�Gi�d�R�49"��~�(|����9!�m i!�����+%�%�����r�	�V�PJR�UU{��6�k�^�r�6��z�gע����j��~�G�G��x��c:a�:�N_����Z��Jd��^NY�g�	H��C��є�M�RX)�y(]8w�Cp�`�ڻh�+�\jm������g%ITG����mF�t,C!����|v�Fy�|a2���54��y�F��[��9D�4��d� #�fN��Rۻ~n�8�ǙF`bxno��HY��'V����O+H��|x���Fʀ�jwWW@tO �h(��fs��Y_�����,�|�<�����\F�����f��;F@xD���Նѣi��F`ҥ1��l&���Q`� -��1�/*�F[�[-@K�D���,<�Z^�N�
����M@�A�M@�(h�ϐ�����(�>be0Cz�>��g
@�k���P`v��w�g(�+��
<�S���A�������|o�}�N#km�ȟ���U���ښN�����-����gr=_�k�Nɞ:t�X[��Bt�_�����~V�l_~�e�1<����;w�`v~�#CZƕ{q����������;��j�h8���4�$���+��:�i���BmQ�p�BCB�������=Ffa2���u�E3����`�[��M�.}�2� Ͱ|����|F��+<_A�L���YO<��_�>r;u��[{[��*E� ��.���WU-,���I|�c���nY':7v6��z���m|���ݸp�9zf|���S����J�&�}�#��YE��ԥ��A���g?��x�?'p���b՘��S���	,�?��.������(.|�y|��߀'��c�u�`m3�L��c�.��/���x��Hv�n!�u�$�H뵣ÚY�K�0(�6�Rm"2��%-�?���p')-(<��[��L����iU(i�3�g"���r}���Fτ��1,���H��'8
����xO��L�����P���� u�n^����R�5���f^��0��*
�����8��i�f��*��a'B.+*��m�Dۥ~��?0(mq�"���ዸv�-�����"���X�a@�^F��6�����z�l���G?��*-e�Y\�y+������ݥ[*_xfqۼ��N�vo��]��R�&���2y�&%�"A)E%��3���B��e�B*n��䞕
G�Q�J��뇃Q[%��3�EQ�e��a�JƱJU�!�/�Eđ���l��]��pVi;�<�"���}��A4)K�C �d��I���/�����b�6�#̦D��a��F�ؽ8x.�#��CȖd
}T�˼Óf�3����B%�{�R�j�̀֡���n_��$.�/��<z�����֚���Ng�P��.�5J��h}��эݝ�:����V|M���j&�k�=1����Hm����*�'�	�$�.��]M,.#r!@uZi$|J��ؙ�idiW:���)�P��"aV��`H	�<����~'v;h^z�6NP��ü����~W�(ꕴ�D}��=ؾ����a/�
���&e��b��-���\���'p:4��Pl�Y_�|7�_�S��p~����oX߸�G�Ѯ屺�P/d����s:p"iց5�vO{��mn� �-h�L�.FH�:�ϿG#F���,�I^'`Jd��:�hy�~��x|>J%c# $��lZ� ��1�O�RtH�}z�q�Hgɧ��P�Xd���� <e��r���_A��E���S2�F/�d ;�����ޞ�cө��IJF~/6�В���]&�4	�l�H�LH�f�d, O��P[���`�*j�%��յ�%��๗j���+�!9��=&15;�uu3�����0#c��O|VK��������R���6��2H ���L����/��?����~ٴޱ�^���Tzl�⸖�-"*m2�[�,^�H}�� <#�������}:�2�/�棚E�'��ӡKiK䵚t��j�.���{(U��tM3���u�x�C�����t��7qb!���z��(�������#
1��u��Џc��"�/8��BAZ�g3]�g��|˘^���^�|��%������'>��I�5���~ϯi�^��O����ʡ\L�O�.L�������l�oa��S0;#��'�$	�z*�&�%���+�,����OT�Tu
��E��_/���sըWt!2�5a�Xlf�1�������!��U�DVQ�M8}d�O���̬M	����:�P ��7��lC}���������h|�9˽G��/�б���?�=l�;�N���P�a!p'(�N �*�z�[m��v�ts�AW"��$��}䪻8<3 �����o���F�X~��!��S)��zg����������;w��Y��A�\@�m��xB��j������8D;[T����F᮴�ￌ��q�k�픸���_�{�Bb�kX~p�ΞT�����R�l�����~�Ԥ}�&څ�rӊ���e�+�wlS.���Amz��+����gne�U�N��(U�>�hC��$����`rExvbZ%��>,^���8}	>����!�ju���X�Z!�L�ٸ>Ӿ&�Rn���ɠ_FԱhs���4�����;1{�:����-��#	H7	\��(��ry�	�>4�c�&I�[&?A�G��{<����`i����G�G��x�&f���Y$뢲m���2d¸ӱ����PX�����01
�-��Q� ���z��4���k��S1�O?�1dV<�ݺ��� �H��/atv�!b�	F�ˌ��Ӂ���o& t�T�bk3��OʧB_ }�V&#f�`(�E�SC�����&���n
��^7#x��w^�ʃ�	���d����V�������;y7v+��̪UѤ��8Вi4�ш7���4ogy��~.����<�%.v�7^��W6���?���cP� W2J��VVd���ֵ����6b�d���,��p(�Z)K�N�(���k�H�L2X���'y� ��KM�%e9�̕���(`T�G<
(;�$`*)�R�x8IFT�S���wJ��ν�:�+`L�>$󶲲�YIy�A/��V ^��0�����
�Wp��,{T�������y�YR�6������!z���s��f�"��dU�A�we-�Ffuu%�H$�׷��ɵe���O���;���KJF.S�%�>���II�F^�z� �8.^|���Cf����pl֯�Ca�y&'����A�d!��j�J©�(�6�����ش�Һ�`d��cV>�
��?�.����/)���@)�e �G�oA�@��sr������M��A+w��uT���k�����4��g~X�C�ܾu��Єp�G����D�~�M
b�06w6�7G��x��a&��cs�[��4%[��UA���Lz���b@W'Hhtt+�M*i���-� &���a��Ə	Ї(1����ݗR<׎���!��y]����Ctt�@dUώdkf�'Q���!؟���k��'���[+��կ�W\��S�>�uk�0�Ӊ�Xj#ȽVHmh0`��:P�ٍ��t"!��d:�~��̙i�MN�%l����C��#�%�܂�<:����W 	�h��o��d�A�����+7�]g�+����:��G��E�C˟~���
sǦ�rg7��^~�Ajp�c<��m�9ޗ�1���9B�����\Py��6m�lѡ�� ��^�0Ao�J�
wS�?��?�o�
�k����T΅�gFk r�5t��!��w;u�v0�d�m��q/:C�0�i���C^H{����v��A"14%�u8x�"m�G���Np-b\G+��4��nHv-��$=��wPˠI.e�ë43چ����B�.i��焲�b����Q��eڕ*ַ��[�z�z���O��s�b�B���ƈhU��׏a��ػUmk}�m�r�-�v�����W���Vˣ��G��x��ͮ��Y����M{�Lq� .����U�N%�����sU:�Ey��k�H����^���r��޷��1'�#�b.o���=2&��|F�^ʅ���'�
��F���p�E�I���0*��gT�����4��gj�ug}Y#t�?��m��N
Ww6n�C«��0� �����Xh�C!v�;t~�h��$6#ہ{�I��L���_�! ��>���p{�2�/ŋ��=�~�~AVm�$�����ڄ,NEz�&&�t�EcZ��%�(4�� ��T�ch8�^yR�ÇѨ74�&�
 �.A�&b�%�����g���%��	P�l������=	X\Yy��L8���� 0���}n��]��QܻwOޡC����a�쐀Kn����2�P,`����e_�Һƒ���+�T��5{뭷�x��^��Dv@�8`���{����<�;�<V�:5׭��|o��n6�I�)ҲlKb$9� ?�� �� F���F`��a��%۲E&�IQ$%�ɞ��Ýǚ�3���[��������Uu����������[���(��00(P&���zv�҅T�"=���w৖�������u�����tQ�4�f�"�����ý����/l����\O
m����M��?�C�������غ��K�@�[��6��ޗ<�O=}���@�����)=��8��P0�.�D��J���5�h8�#q�|�2�	��U���F��sY>k���Lz�,�i�F�mΌ�zU�5�x��ǽtM���r�%i�l�ğ���a�����&�IL��\�M�O%1��)PD��آ1v���HL�R.#� v�?��Ic���s�}��p�O\$�H�������A	�gp��}���S��C�ڶ�d�pm>w�եAC�s�\5�%�{{	
�]��R��f�1S�[�Z��ΰ��MnӪ��^<����#6�Ā���E�V�^���em7E�!�TU~��#5;m��D���������@rވ^��Շ{���Y��N���&�CSI/�̀kE�
#I���8��.	G��^�z��>�%�������;o?�2�e�@K�Bc�i��@A~C�u,|.��77�%9�6ڛ^��QG�<Ak�p��&ǯ�˾�кu	�B�>�����V�������NF��k4��HO��{�c�m��U'(G&p��&*�M�9�A�Z�B�;����4��Ln��h�F�©�-�[�^�@,��� ��A;i�.�cQ�3�Sq �`S�^"5��}��%13����.�wߪȷ�r��_���c/S�&�P8�2�;i����K3��>h�6+4��|W������Ѡ{@��yl��/��x�ޘ	��F���Ò����~���� �|�6�<s�����'N^����0����p��yc�7zp�^�4T�t��)�y�ln���k��B��VE�3�[����h���x|�
Ǘ�mgWE&N����I�,��R7�ִ�ବ����b����<�C
��}��ǈP��on��/��ڋ/�ko�_�W�g�����hE�L2��;��/��@����������up����O����}n�a
�A����w��j���
Or�w��8�`����xC��G��9
�N]��>���S����~����B�A\.A�C�ԅk�ϣ1�pǋ}��ԔA*�ΰ��;�p��I��?�����PP��?�Z�)��ͯ���hYa����gx���w�?���o�sR�<f^o��%j�W��r۔k%p����r����w�ӌs
�ĩ���t�ʕ"����y	%X��Ԕ����_! <0 x���/r5�#O��(O����������G� ������ ա@^ʽ�����bU[�_�8Qc(��N�!�)%w�`S3]_�חƩ������ӧ�*@)�'��Q%��p$ �-��e��T���;�G��9��X<��������'?�Х�*���c8���~�C�y�r;z5���->�]<�̳x������q���'�ҦB����v{E@�3~J�qX\�U�>8�J�~F�4�p�n;���fQ��T$9=�|&/�w�ZʠL���'iP�po��p
f�j������S}�!�_�j�`É��98G\4����UC�<���q���8ߣ�t�'����`i>��'	��������͝¡���ޛs�'ￍ��P��	�z�]vo��F�ѤpzEvN���eN�T6��#�SO���AԠ,!a�p$���	�2h���vT5��\y������L;B�G|�0��u���+���{Q�A�9�,���kƈ)��W��?x�k�`'�B��Hl�d�
f\��s�۪
�Z�E'P�W��s�6���ݼ���m�ӽ��ű�Qe�r�*�^�*�k�����a�hܵQ�$�.[���]-�ȸ��hUZ��ڶ^��ȸ��W��%�(`-%={��~��~�C�pO�f���o��kϾ������1�V�=G=72�u�j*ޠ\)U��!!s,E�̸/���-2����Ǩ���~�
�*GVm5�]��n��珣FY�`QO�(��J�:b�	��GM�dK��}��@��y��9Qʨ����O��[e{��4"��DGսN�uL�(�h�[Xۊ�Ʃ{cF�yb��L�q:4dOb?W������������+൯}��������!������/~�K�.µr�-��k/࣏�����«/?M=�"���iM��*�m��4ƕΏ��Ǘ?�d�qW-q��x�hR@��^n�4� �/�0?C�L������V���)�>�!��Ź�el����ӳ�}�R(���2>#�:��'��šH�i�6:T}
n�< �ɻ�ݘ^\@�@*5M 2�FK�5�8{���P���y�~LN����8���q|��;��zGh�q�-a<>�`�����~�ۿ�xz��8��uRA8LX�P��ÇH�����V�yP���@���ME=� nz{x���w�O˿�G���^��߲^�y���m�r߽{�
S�rE�H�/Dg "k+�����H\�&1돛NO��s~�a�1fM�LQ�t���B�*r��"vm	��Ü���0�9w�� a�
Y.	�q�ƈ��o�wU1�"���GN���@�G����}��U��ĉ+�-`��[8�O^Qy	�ԤH���H�]|~*�\6oc�N�X��Z˩{�>��������J^8��Bݪ����8-J�9,W+��|h	���+Fﱹ�iO>�$��&��S���P/�o4��-8��B`]�������'�?ϝ�!E �ҋ�X(Y�!O��k݈�WGnܸ��|�;���u<�y�� �������b�`�F�����BM�Y>C,��R���7P��h4n��&Q<z�Xjݺ�o��>�x��"&��ko��3D�⩫�Q��/-��l�Y�>��D���t(����L�˴�"����9���79�(I�-a��ÃC$�3|��\�׵'��n��_�k���7,5�Yo!���cPS�N��;
���5�2@.����jt�y&��Yvg�o}̵��Mq���-R�7��Aӊ=����k�ݼ��I�`.���Uyɍ���X{�,�_�ޖu�p9�fL��`��bznw>��|�8����M�)y�����>���T�
�[���L4,�Q(�Ъ8̮`���a��$�ܺG�6$�R�sʕv��(�7F�	H������uAYV�U��]x��M�u���b>d��c��!�a��ñ�+���9���(?BHϥQ���/�����+3jM���`Ǘ�8�9-齞)����y�	��,��$hFp�[HMN��絆j���Ƿ���B�㶝C�����P�۾4G�5����p��(�����u\=�gX:u��<\�k>m�>�шk��uDá����d~ղ��W8�qM������W��<{.��ZC�^�������V5L$j�5�͔�ഖs�ϵ���RDo���?J�[�~ �=yw��)�&�'W�r����x�ݛ��zz�g���Cs;���u�'Or���X�ajb�2xрt�Z�V̡�9'���=F���_�����c�L�گZ%V_�
�b��V�e*��?�̼C�)yp������ S�0]uz�uk:�JF�ž�>1���q:��~�,7������U,"Z5X�M$Q�vPn�iY�x�iμ%�L$E�РU_�����B1���S!j�'�p+�(�K(��x��s����M&�r�x�DR<��&��m�
�hŶ[=���:��3F�w������6�wQ�搡 ��������'����w	*v�(/G�ͣ�<0�у,�O^&�}�Y{�X' ZY^�n%�f��.,��R�8˹S~�A^42��~�o��#�i�ɳ��T*���+o�c��w�TQ.�r��(���˗͒`����>c���/i��W�\��ￏ+W/Y��>w����\�����=��4O-*��
۬���y�z=G.�1Ъ9�u����S2a}DK#����4��6G� �WR� ���֜�����8O�:���Gڇ�s�3��&�,Ϟx%�J��������{�<���*ߛ���v���i���_� �:�E"��T;�T<9����e}!�$.�XW������l%ȠB*�|N�?<$X�� P������&�+MDO^���_}���Ϳ�Š�F���g!B�5"@i�7T��!.�/<�Gwo����>w�*+�i̤gy�,��!j�Ж�<W�d�����j�3!�8  ��IDAT�n�p���|�%ܾ� ��_�����A�k^�0��&�ua�fkX>��g��:(6׷	����9�q��m#NOL���f��c��!�-����#8����?sr��ۏ���x������wP��Sy���
��[�ЁR��Oυd4�Q��峽q��X�(�Z��j9��y	ԋ(�s4 K���(��4�4	l��q�I�˄�5�f���cw�!Μ>�[�?6��6��$�Z�c��$ț��2T�f8�p��ȥ�=�x����g�q�*de���=�(�]vz��hWzF���0���^���&<�^�O������(���у�����Q���"D�0Eâ�������m*4r�i�<�ڰ\^�'�u�3i,��>S�{,l�y�s`D΍�Z�90��4�����m?u�u��/�dX+U#�}�7 ���])�UU��sW���ak7�Z1�u:�==�(5{�,�mʚ�@9�-u=&���R�I���{u!S�[J����C�:�`�r��C�-��v�;5�s>U=�3����������p_&17/���u������8~����i� ���R��X��9�����/'X�YkՅ��i!޷4�!ׁ�^���t�>���\����������:iKq�ךۈj���������rSQ�oa��
^��W��'�������Ut����,`k��*�x>n�A����cmcs�3�Sȍ�5n�������S�NM�-~��E)`�z1�<�v���M�� �RH���z��"p�7"(���C�/sz���CFOZ�C'�!1�-�By�~��˟�BesH+`�����z$($ ���)9F?AY�\��G���S�pri��y�{���7~�7l����u*�JT&>0�C��ze�V�Z7�����I�2��c���!��P��Ύ�b�[X^-]WU��慌�0�H�=��ӈƓ�&յ��ax��e+TQ�������/P�q^�p���}S���q˽g�}�@��5��m�do|�F�>��
��ʉ�2�<M��8?�P� ���>'o�B@�=��D<��d�B�g�
Չ�{h�a^��	`��Dca�;�Noy��F�I�df���s�7V!v���U��/?��@�s��n�oX�D�VEf��a��R�z'�*lo����+_y��.��?�	�z�)LN�"H�������MXщ��s/=ר�ro��E��K|N��~���	��UAO�òN\�������\�C�3��T3�Q�*&���N\l��.����^�P${"9��ys��<���eV',�w�>�q$c�x�ױ�x����)��]=ű}�?v�>*#}�<�� �#��6�e)��ݛ?���7��?�����O�3&F~��ˢ�J�ǴC|͙�Gx��'13{�ψ��`���H����g'&�T��6��8G��ǟݶv��p ^#yW[���T Y�b�wV�N���T��ڛ�)j�`eK��@�ko{o���/����r"5ǽ�A�ݡq@}�B� �v����u��o���})79�F�z�Z���|y���=�m�!�2c�_8~���.�4l>��b:5�w��z]7/�;8���O�>�E���z�˙���O4�(v\F $�D�F��kd�i��Xںǽ��\�;��)�2���5�<ڴ����k��g���}�qך%dr�ku��5|��[���������:
�F������&'��ũ�≸�n�s�.��+��nl�Iq��R��>P)�ڂFX�,Qf��{gD����Z>�%QE��Fh��\�\��CH�y�^G�*�?G �Y�R��-�����w����0���FK�j5��Z-�c�w���]5�]��ns�3������G���wjD�~JE�'2����K�����?��C\���|�eꍔ��-�4�� ��2~�o�����ל��.p���qR�e���)�e�
��~v�c��ǯt|)P����1ǜ��<T�m�Y
�X�T��7�+������vV7�я����{[Z~㢍�l�h�F�BZ�LhyR1��#���Jt�F�0Z{�b��|���/{FF�[�P�Q0��#�j@3
�û��y�FŁ��8�T<���Ѩu��sA���l%����-�S'���(����|Ԯ'��&U�Ҡ�FA@+�C�4j���KѢ��+/���"����W<����p�8�^�{ￍH0����[����G��:<zH!}��d���>VHsnf���J���[�s�-�gP�M�O^/AY��t��+W�[AI�X��MLL۽U�"��s�=�����b�����מ��{H��Ơ|C]C���3�=w�I��[�so߾iy��䢊^��s��}�/���8�(��\���~��6'/�������)*=�����=���й�c̲o#���Ĕ�]s�uڢ`�"0��������i�pgw�*�UP���V��h_ҩ)��m�����X���y}�J&ply	�߃�3.�x��繢=lo�X^�+�	""t]8}�%�omr^�|�}f"c����-s���>�õ-�	�f�	H�|G�o߸���3������l��ٹ��W��*���"v�|�)z]�u��V�w�P�e��h�.���_D�T�*�Ҩ�`s�.�!��;��#Ɖ����BWr@m��ܧ���$�ı%,��"Кå�O�����3޶ݝ$�/�;N�����5*�W1�BG4>�z�>|��k�T����A��EΝ+'�"5�����k���������dr����N��uaj:j�8�);���J�����{d8ĢIl>Z���y��������� �&פ��}��O?��,EC��6��*F���)�D�(���/?�Gйx�I�
����O�����c2���O�8"<�qi�o�i�)Y����E���qsr�Թ��#(6M��vO$.^���E��Yy�?����ϙ���D$�l�k\�5��X,	OP�*T��v���}�<5��U�`(��ƽ{��:�\�:p�Qʹ0"HKO%P Чل���	N�_�W����ڝ�3p�z�f���E= Â+]�~*���ݪԭ@H�>��T�6�.h ֱ�p
�ܘ�0����B����5��yH3�;�'�nL�
�C�����RC� ���Q\�]%VU���yD#adw(��s^�4"���!��E?��;����:{y04N�6�N�2����w��^����A7oܣL{Ͻ�-+����5�����0�i�U꤯�7�C��.^^A�LÅ�q���������(i�x|<>~��K�B�7)�֘�����Zr���z�uGF] R�!k�u��9������D%Q����>��gLKT&q.�	�n�:q�D*�y���R%E�ۦ����Om�Z��`��ȩ˸���E\�[y�&7j���
"���f��Z��/��ψ���m���s�y}�	���l�y,�kg��S�)��)[Q{�9"���&��Y���_x�r��~��Ο?� ��v����G��ؘ�P���y�ԇW���$�66�/�~v|��N`\J�W����� ����m��)���A�Y_�?�}�;,�,0�
�+����@�@�<�G��K��[o��Y�Y%��{}����{'޸�]������u�)��U&���B���%��zFԪ�Zi�k�G%(�)/��&Ч�DU�" %�l]J��c���Qy�w�GTXX�.�1E��Z��������q(Y���<�G��5�N?��6?�}l��g���^�g�|l�W/��;wnYQ�`P#0����~� )�kO�����G��0�6F�H�����e�!W�{͍f����SW���'XlR�����(QY�!�YDr�`J�w9�S���T�%L�Sx�xĿŬ�V�Z@��9{|ۛ�H&���Z��fQ?�#B ��c��&\?w6p��g�E�@��Gr:����'��ej>W�k��*��Z	v�{�4����V��it�Y���%�[�������m�+O��528w-�g���W���^xuL��w`��E��z��z1o]�(D�fg��z,j�$J`"7/���<�J�)D	l��8*��¼��
�]Mb�sD� �~��G����_z�Fk�\�<s
�N.������j"�3�%ivU��u^�:e���yܼ�!��"��9ۏi����k���}U'��Qլ��m��x��,2�A���G���r�0�[���˩\7�_֌��ýX��(+c�;J��~����6FOt(ێ�+����R��j���[jj�r։�>x��nޣ?�����=�F� p�{r�����F�����b2��T���C��v�^��|d�����z����U�pv)�.^���+u�5fѢZ]��H�pW!M����bK��%|\����F�s��֦���UZC������	r�['���n	��9���Ġ�ȴ(����u�	,,������h[JS�;.�[��Y*�����\E(��(h�R���7��mTۮq�\8��E�D0��x�vNV��~ny[;�{��?���:����eS�D`]F9�.>=KRK���y�O����s�q����_
vnG��i!z<	�-.H�YL����Ԋ'?�X�Rf��7F�o����8��
���"fs�1��[9Lm�BAZXU
��ȎV�Z)�G�c���C1�z��θ���㰨�}P~�ZE1���CPX��r��HG�N-DZ��F]%=7�'������7D!Z�S�����A^��J�&���J�S���[����ƣGo�1hS�-�Y*�GH��}f�ϜDp2N[��;7-�* �J�BavTZ��0%7K`&С��H�ԩ���g�����N��:s�sY�cS�V�L��7�|�@���9��ޝ��~'Zy�2�GP���lL�`�7I�:���h�;������_�J�����f�l�s�k�~�
]|*�_�"p��鳺��U�&���u=)k���n&z�|~��%�vTa<���Au>7t:R��7�
o�l}A��б �ޝ�R!l�Y!!)=��%�~��
Tf�MAˋP(����}��Ξ;mϡ.'�D��/�������Shr�lng����ď�Db����]9k�"�}��W�JRi�y��V5�<b�w�S�՟}��]�1��rq�
w���U�}!�(in6�v�c8�(/x`��"�Q�^��0�����E3�����.�M�ް�آU
Q��h�����˃2��5s��Y7ϱ���T��T���Y[��n>@�U-��ͫ������
xf"��Qq��lz����{vrʈ��>��L�r�r���UoXzE�TF,5���!eɈ p5ʝ)�Wo8��7�t�PQ�/�~��G�-+��QU��G��o[�7��|�`b�w��Ň���(d�X{�&�QC=�G��[�7D�@�T�Y�[��ec� ��$b� R3S!|���q���Q�� ���6�'ɷP� ��Ba�ay���$
�<׈B�~��=�9�[+���^J���%��B�k�=j���;N��"0۷�ȋg/�Ro��ޓWqd���a��Y���=�� a1ߍ#`�5Lн0�}���҉��T���D�z	s��W����g��"���zݢn�a�H����qOH�T���e-}4�.ʏF.
�����J��szP�)Ӻ\�!�jUL�)+�
E�bR�;����	�t6���i��p|.�A�E0�B�W���h��\�Q}j�PE��%p�3*����E���5�'*}G^J1+���ۏ�7a{^t[�|/��@}�ڦ+���!�	�#�	���ZQ��&�-��.��rwt�|��q7Z�q�yo�h�a�x|<>~����pC��=��ATi9��7�%��c2}��d�$ܦrp;���B�񅕅���L�u�
#�ť9#n�� ~���%��j+T�Xʼw�f.Bm��gd���,}�N�g������7�X�\���)��;���
|."��vh�)?�U��Qo�V!�mZ��T��3�(f+.Kp5he�S�w'���������O���@��G�2��% �r�Ϝ101;���l���O��Q+�o�3����8IYBD���X���	�@��/ �q�=z6��D2i�.^0�6�����������(��n�-�+��{]"C�5��r/���U�
�(ԫ�$�����y�'�
=^x�����P��%�/	JU��cy��=�Q��[ȼ���ʋX��(R�	0���@��)�yn�V�0��wDT��Sդ����A���z�2��g����޻3��ܸ��ԩS��|*Q�(��C��I�X��޽����]�r�n�B�ƍ���?�1~�w�c@��?�!�=����`�;��P ����+I��B'Q]�t��ǈww���֞J� �$(S�]�s��������8~�8�\���y��w��*�)>_L㖁����7�:�נ+j� Z�ݶ��X91�[����W/pϠ�����Y�	�]���5Ф��������Ki�]����ߵ.+�a��t`\�6�`��-��<f�g���b��X%0_Z������=�p�Nǁ��>�?����p��!`�9}�YxBcoI��f26��!�`�����x�w�ݫb��;�K-�����7,��Qo������0>�d3(�!��UZn$����:�V(C�7�߳�í��72�J��յu�:	z;�s���d\$�F�U"�V拢a�`Ə�'�}�#^��>��k�����o�FM7�3u�\NZy�gJB�h&s��(��\_n�c�Q�����pb�d��޾���~P��]���
������f�����=p�{���M8<x��BD� �jmʯ�7����u���Z]���9<������?1� ��1E�o�Ӏ���\]��'�C���6�b��b#���:��}e�m��)��[����d���P%	������Z�h�H�����Z�A�w�H{���k�)���#����8�pk�[\?����&݁�����k9������kN��m���l���L��F���4���z�kV�)o[KJ94���;�&6�K��;8�<Kq��;�nqV��<c|����ɸ��T9����	-/<�+|||��ˁB���"�����U�O�^�RT,LʹF!��|	�Dl�ڶ���s[�������~��y��u
��Y�	��ƃ�Di�S�q5Z]�fSF���DQ��[m��
����P�)!Z�T�x
��%�U0�
P;�nr��*�F�O|>�u��S *t����eU7vp��O̜��>���%����-�|��?�G!]�bj~�p���SO^������H7X��)|+_Q�D����j>�h|N� /�Q�6)Z��Z��Z�
��k�A�����+o�>�/][�ɛU��?oɤ��-�N)�(@�)�#`{��U�Y�7O��:X���Z9���[&�* ����d��\�ɛ�P������ ��u?�{D����Z�����)B,���-�^��pz�.(�����X7�q(�R�=]C_zv���H��M�]���g��n�;�{oj5ߺ��6�aT���U�.`�Ǥy@�7��yM�N�B>�)-B��j���e����M��������u\}�U����Wb�3Mu*����������q�����7������������2�ND��^������,b�����{�2D�����\7T�wCd&��ÿ������P-W��<����������	�h��`;u�Z���<�I|��g	p�n�:�nO=qW�\�6��B��e�m�}ƽ����@�w�ӿ��מ3�og���f�ʋO��_�����wx��OX��v�<������y��w��n���r8I�CH:}!��i��Ѥ��,�P'�_��?���6����ȖCϾ�U\���
r:��<�Z� ۅG4zUD2u�O�a�Vg����{�$��"���Y<:����Yʉ�\�~Ϟ��+_�����B�'/���]��Zu��Iښ-8��|�bERS�|��c���#�������'�����o�|�^'�cΊ�"�$(��Ny�^�5;h�){4.R�#�=,�ߠ1ܺ���+����q��r��$�)�{Ϡ������r0�
�G�&��5>��DM�;�3�R�d'�y����|�<Α�	Uԫ�~��,��O&��V�'�AcX4`� ���a��ت#�#��Z<���;�}ei����6��׌x7��P��M}Z�oE 3��5�1��z4Kf{C��>F������ ��G�)~���
�ԕ�#��u����'�������5
��|7n�|I���W�
��A�:]����o=�j����Ǘ�)�u*�9�bj�f��@���B(L�Б�\��Ń�w(4�hS�9�*.�9��*hm�����Kq{�ڊ K%'޲~�cd�w�~�1e a
+1�K�IpF��]�A��=�DK�W�X�WA�@~Z�#51wZN��+2TO�J`d}{e����>h7&<�����#���@еy��K�}������g�ǩhi�&�TrE�@�ĕS����;����Bp���c�	��U^�x؎:�(�:&l;�7�;�*}��!�|G�Uy��x�{G������ӡ\)kg��m[���ƪU���u����az������\�B��v)�N�B�>vP���� ������,ʱ�8$DE��0�@��XV�Z�8�ҽ ��;
EQ��z�9E�����<Jy	u?}^@N� �,n1��qqH��r���:�����{Q��ĉq�Uf�Ba����7=�0�Q�(LX�g��4X��{@Pu�`[;�c��O�\�?�[�X2�l)g���I%�N@��?ķ����0����
�Di����\����B���/�{�w�n���ѿ �O>�!�>��n��6����;��9{ߊJ\I��"|����T��~,̈��-�:��^��*�;�B��ѻy������
������Ԅ�G� BW��#<sr;�h�����^�72IH���3������ͻ����S���A���$Ƿűp�'S�ȣ���+�-���51���v������0�JmAA��cy�2��"{�ܳ��e��ާ�����*�]\��B�{��J�s!�+_D��D*��W��6^��>��-ܻ�� &����r������Dl�j	���rbDr�sb*|�!eA$6��_x��f��h�^�2�$ ��_�:�ch�H"��(���� "��v� ��
�(���)�9�|�
Ο�j�У�&������r.�l�~._��$GΎQ���s=ex+/Ǆ��1�/S~͓8 ���T�p4Ѡ&hҾRITQ�(�P���m�A������ȡ���G	�C��>A�l7�f�U�w����E��.��+�ZA���Q���i�W�2��� ��z�xy�{��
cL�����U)������
��!8}ER�i.��]L��x��j�@#M��Q��D�.�j�
���sա��*!�x�<��h�c�o���L�WP=��B���8�$���Q��߽Nc[��ΧZ�{;D��i��{��*��#ox4p8��h_����&~Y�#�$WI��H ����kH�8	�f	�FV������d�x�\���mV��T�����+��x�`'O-R��z=AKwb�SY��6����p���J�]b�W�6Uz�c�b��59�Q��V"�O9m���Î(���Z<oHp�H���(ҲLFpwk���e�:(@���|�>���9l����j�e��~��vn�`Qo� �X�d�>|.*��Ԭy�d�8���x:�8YhS�@j+ǱU$���ڽq^�<�F��9��@������@�<T�� �_��_X�C��uv.Ñ��D�g��!a����uh��Α�QӵԎB����g�<��_��#�@Q,5���q#����,������P���w�Q�����yQ��;) �{i��5�G�Z�Ty�J)е��Խ�}̡�/��:O�S���ĳ��)�뮯mY�f*==������dye�m�q3 ����:pD�4�����Bv}�	^}�+6�O�����c��o}�B�����ǫ��f ����`-�Ç�ޢrN��է�#HT���Y�~���c贫|�&��:܋�����o�̉㖯�	Ю��F�a�W'0(c"�"����-8�#ܹ{��h�L�V��Ƨ����x�x{��MxK;XHN��?@R���`s���<j���,��S'(��ԹK��������F(�$`���;��-`~f�J/���()���hً���5tzU��L��$	,��B��&\�����Y���EP�[��ĈcXJ#0<�v��氂!�C�7��<��D�N�v	V0�D	�'�|O\{�Z�5���ZqF����9��4�����3�"�����H�����r��̉a� ���E�y��ffͨ��'�Ü���>����~��G�q�����;��Fp�4�o�ܙex)w
�v�e�.bz���{o�����Kd�������,Sn��ǳ2��A�d��I�RuX�����������w\�&��YTW1T�8�����Rζoܕ���Eh�[�C�h�r"h_ƣ!��Dbze��r�
����k^B�E��ې�@�ݢ�꨺!�C�f
q]�h�����
����W��XbW�	�s8srg�ˈz�X�@�z� XEj�J��8CC�G����0�����R��F�&:�Ѹ/�B�����\'��}�H�6��+�Zg2�b����G-_F�����"�mZ���n��+i����������l����%������+_
�F�рZM�<��`_�.�=3K�XA�@�<& ܵ⎑� �ō���f�A
�ny_���S�1Z�[HP(�	r$|>*�<<����rP���ϐJI��33s��M#n����km�Sxe�vX8NBW�M�zGjr�M]Sk)Z��a�V9��FuZ����"O�a��F i7[����_�]4j*p��H�������Z�X��1���`���A��������Z vh��:PmE�������C�A
m� ���R%��č��L���bY��0���¼��|L����ZR�+Х����F�<�Jp�S��:�l�1�L��?4�l@K�'���՝���;fD�SR2Z3�s��������5���y4"��\��<
-�����~��u�x�}$�7�-]��z���2/����4Σ*d{v��]㵬ߩCL��vLS3a�]�Y���S�>ok�q	xJؗ+C����Y�Z�!T�y����j36��4�3��vbv� �r�:���8��|�Vü�'O��W��rc�����|7��4� T85�O=��s�p��Yll����?�$�~��m,���heַ�6�C�F�Z���79fyӮ��}��g	҆����]��ۆ��Z��|�+ �g�Q��W�2��B֯y�&z-D����xqX���}�n��1�����*���)��9,,�@�YB���"�ñs���r߽�z'�׾��)��aͽ��g���xwc��u��5�����6�8�q�-�`*}���C�/����l�܃�W(�ֶ�L \�q��$	��h�O�G��DX���#t�����x�̦&htR�JX{��R�S� ʹ��h�:���?A�!8ߩ�E���ɵ�}x�f�Rgf���h��-,̢Q/ t1h��F�|�{o��<��`"�\��ȗ&��K�����Q�;Do胻����fN�q�A̟:���?�;�{�S&��&`Q�AM�VAz�� �u�QA� ��so�&!��v���ƅ����7�����'����:
��A�"D.b�!|SQK�֊H����۫�8V��/�^ߢ��&���Ho��8��0��'d`x�
r?�ᛘB�������Pp�C`�A��f5�|�����u��h�����gރ��v� �\��ZU�F^�do��~�F�
\�nU�SN����(B5r� ]t5�ߣ\���k����p��W037M=y��y�.� C}�NqbȖ��(^]���c�FV�F��:Mi&��4�7p�t���P�,��"�P0������+_
��K���P��Z��AuZ7>kYW.e��[�lSӓ�6,/$J�K��F���.\8V��im�K.u둧Q4��G��k��Z�r�\T F ��v�:�=R�٧��N*L�Uՙ�����x���K�Q��}ρ`z2���C"�B��Z��^ ��+�~���AØ�̃�N�j4���YT�yLS��(�M�!�p�lt͊��Ѯ���w���OP5�Byǒ�)�B	��s%�p�>���R���.�JZ�<��P��D�kԚ�/>�Vj�k�X�{�g�z�hm����PO`:��'���~���s�Z�P����z4N]G�>����WO��(Q�|�+�C�UdK�(�Q��=�]�f-�4G��. ,Pjt��-����K=�u�q^и�E ���GU�:_���a���>�{D�u7��#�B�_�jb.]���t�Ƥw��|�:�,o��I�f��c���n��%*eO ��{ڽ�>v�o������ۺ��z�k�gҏ�.���m<Z�w����"q�P/<��0��@D��gO����x����k8�p��;�'._�t:���uܼ�s{�Q�j�4���^�^w��n��Wo�yu
���@��7��s�R�<\�3?��c'(&���ϱ���S��5��_��IL�&p�D��#l����;��y�6�)e��:�y� ��`�p��c�����cv~fL�3��o��T�|'#
����X>������?����H�G
3��9I�8�.����c�O.o%Ux��x�� �8���mI#��Fn跜�N��Xh�y���W. �s�V�������0���ٿ��qF�sl�4J�;|^ �wtp�����VɈ�u��2���;��o��<]��M�f�	��}�	���$a?��/�������y_����E��	@A�Ǭ���a4r��}��R|�3|;;wP.摠�[羙���lӃui�x�G��qp5[��g}�Y�&#��(J�CΕ�
q��\OZ�n���5��>Q�uT5��鲂�Awd�b��|/��4j�}_�	�-a��^�ǖ,߼R�А���}&�/Ӡ�T"�k��5xM���M������KX�9oȁ��C�U,�M [m�#) ,��gц>פ%��Ɔ����{t�;	4�|W�-*<��;���qS�֖O�0�k��q6�G7��/^E�t�����Ez>���{\9�O7�F�S�%��F�������+_
�Nw;�C)f�U�:��Ր�'O�8MK1�-�*ԙ3�T�y��ݡe89�x�x����(�똝J�pw��*F�an:EK/O���;��h_\���[}P;�B��h�7p�K�Bݩ��Jw�sK�FG#Z�N%8{<���B�29��p{b��0u�����'����=�BN�L	��^�l���`�wy='w� ���yE9	��g���Ӱv�1��/��+R`���z�����,��($*O����� =��e���������B��o���3�X��ч�{��9k:W^/y�O�7����ј�����g� � �@�r�t	�db��{����TE<}��(����~
��磼F]G=��iܹ{����w=��gG���ޥ��)���
�j���<�ks^��\�*/R�觞�f�I�[ƀ �ŋ�����ٽ�ƥ
c��� c��
I��������#�/%ٳ�=*|v��ic*�뗿���t}��(V�A�X��Uk�B)uc9���]�a���ķ��7��|�K��7���͝������7�/��U��ˍ��]a*�z�<�+0��a���u��ܺ�j���U��gq��Y8z>��]t�E^?�
�nB� �! я�>e����&$���by����Qm����$����{Y\�t�ʳcm17��,"�Yn�.N���$������vsv�8C�Zn50��%(Q�5L4��y� �AE=�����|d�W��
��W*eʗ-�2�Uvq���F}��%h[�hzpPT�,��W/?�ɓ���=`�A���}��<��h�9�x�"�}��%��nKw� 8��Tb�Ss���w�ٹ�g�x���QW.�"����7��{,�# (�������i ����Wq�_Ż���rn;�2<N���r�a4&2Bu�p&���z�)��0�����:����U������<ȩ��C�b��t|�(�i�/�V�1=�H��e�).kE��{��'(��#7�ɰC� �d���N���w����TY{J��uW!�s��0B�ѷ�5I������E�FbHr��r�2�h|�a�Ys���~D5��$����Z���^�T',}����
�"@N�g6���O����8~a��*�o�gnqf)��ǩw��	7����W�3�B��0�6���"���z�
�#������A�"�_k�n��`��X��;o�^}��3)�"���zg�x�,u��>���*~�?���6֯�T���'�h�V�n1�^���ݑ���`���ǯp|)PXQG�^�%/�r�$�D�R*挳0�#�bk�b^����DNM�̫"��V��[�oS�{�Z,��T��[Fz&��Հ[6�}��e�V��#k)����9���;j5'��q��G��vqTf��RT�?N�W��B��d��7��LRV��i����[�bX(�Yw`2>�[��ý���v��y����������Ū��>
��+��#x��M�gU�Q��'o�B���q���V��U> ���JaH��	
d]/L�"�#��<v�����}G���P�@�>/��'�Q�>/O� ��qT5,��C9��������h��%� ��S�Nޭ#�l�]ͅƤ����U��~֗����D@J ٪;�/~���~��.X�����#���M�՘.֜ȣ�s�
����;�Ж'�h���!>?�e�U+��<���	+�K����iT�*b�R˯�<�T���j�Y�8�S3�##���Ɯ�"#W�À�9Kp��;��������%��\�d��>6�ױ�>eK"����*�WWa�u�k+<��4{���N�����g4�v����?@�ҡ�v�N��.�&�k��Jr�@�]:���u�;q�Wqc��@��J9�{w>Ejҍ��.r	^�H|�R%���^d���T��r�=�^a�O^�{ZC��$�^!�"�����<rh��9�Y^7H�6h 6��K��;����;fؕKLNM�P�� gO�'p����,��M�&�y��k_ã)�"�p�%�A\͚�n�Fa8��u��3�?j��﯐��Ǳ����� �T�o���bn~��>�?���ͽ��$��ѩ��"N���zAg �r� �sr�h���ʫ���Ͽ��9|�[���wh�UQj-ҸS^�r�¡���#p��yWN=�5��R�M�p�n���]s�k��ύy��>��ҩ�U�z��ArF�[s8N��Y�������CU*E���`��շ<Mذ3�^�D9X�2�Z��*�E����8�\���`8s��M9-�����`$��1�r��g(u���Dgt�n�a�-Q��䬮m��2�?a��~��PPd�+4r?<a# /Ґ��)t��'�������r�{�.��lc@īT#G�m��\�n��6�=�i��W5Wन�C)J�j�Cmʕ?/��b��V- =7A#����;8�r��$�?��O>
ᅗ�ܣ��z�թ�hLn��O~��frH�_���N���q�8����p��$�T��x|�
Ǘ�}��`v;Z���FI�uR~����sQ�(��!�SX�,,�o�Jμ$֝C<v>����U*�I����f�Qe���A���%'�>��e�*�F[�It5�qۮ^�<��/�V�e������A}[�sc�8.\��UV'P�R����sk���U������� +�Z��f̊u�{HPa���Z�ݻ�ѥB����X�U��Y�e��n��C�N�����L�si �:-�R�r�,Yy84 �cw{A� ��eA.j���L�*�<�����yvt��# �.$H[��˙�E�F��s�s9??k��:_�	�#�i�)����f��<^�^�{�f�T��&`5NY���s����:�DksT����Qٺ�?�E�M`v�W�����G���imʸq㖍E��~/�� ��@s�9y��r�������r�ܹmZ���޳�]z�x<9��������i�j��R�eksvv�<�z�~�kH��r���W�e>��[_H7c��G��/���W���u%�N������ʩs��٤�L�fȑDq$b,ɴ`����a �0� `x�����F��2%R��f����V�9��s>^k��?7_�o���s���߷����{�C~���ֲ�a�W�:���j۵��˿l�*����v���)`��}�=Hw��ŧp�>��x��������_x��<N����~m�s�¥K�����Y,�����N"^q�2h�7�D�k��s_BblK����vS���?����?�n�j��l��h��'�TN8ћ#����'�19Gj��tt��;h�����I��ww{�~N�Z?���}���G^�I�e��|N�x�C>���*�S�L*0����p��$p���"���/�?�A9{�F�e���� �x��l��t�籹������0:7�qf.�����I�B]���N͟F� ���"R#��s>��6�����Ӧ���bm��s��#:����`ԉ��:N�;_ׇ�����6����$�I��k��G���򸰼r�@�C�3�=>ci7�>�:AJ�P�&�T�h2|A^��	#10����ʏQ.��|��_�tʶ�c�~\>�n�x��2Ņ�ƙR�
�P��J@GMQ�`�G�����a\��Щ>�X���R
�`�#�x��7��,XR6����}��.���	�BE�'�`@�G�����\����}\�B�Z_���=�EP"`��˦���l��U�m�n��g-�Sqb4>n�����t��D_�ٙ�\����v>e�/#1wY����1�������h���}�B�[_Pb�'7l�6V��#"��=�!<Z�D�`#���]���2�O]���3�w�*n_�C?t	M��X��5xhr����X�@��7��K\�4�w�2��P]�*CQM���Ģ�"��_��|<�<�z��d���pA���è3a�y*��������/��ne�@�N��FSF��0��`� ����h���z͠_�ƿ��`ˌ���\ �֒���ma���p� t۟vǪ��S��~�@#�I��E���`qi��<�g�yºs�<�,,���A6M�rh,�U:�1���Dj5ܿ��1<��S��Ny�κd��Eĭ앶Tk"8Q&id�8�iSe��q�k�R[ �+n�rղMG��G��F]�)zh[t�c�˪��2i��e����@Dj��3j5�X��ܓ�3��O5�u|
�Z�vjnQ�K�WN�k����P�%m[��~P�R K+[���e���Pe�T���*�g�G<����Ӭ�P��kZ�P�֖��_`�HaE��v���o@X����o�Q
D.-�d����j��e�4��w�9��9��;RK�����}��8��%<X\2�/:"q�����̤���\��OXl��Ïn�- ŵ ���1�g���pwǶ����<���2~�����tOZ���y�zOҡ��?�!^�U�9�������92�7p�g������;�}�����;t|{��8���j��k��4���W��p���xh������!�q�_��j#�?�ܾy[����ۘ��C�q@P���ٴ:�&��"���G~�����w�G���͝4�}��>������q:GigqW�~�_���b��ݷ?B 8�v�G7�y2�~�0
5m񷑈bw�$<�pH��=��%ژNGܛU�Y�� ����c{M[�O�%�t].�kx�p�A���/��q����/�����|�k����������cXy�OЏGk+�����L?�^)e(	�O%��{u�ԅy�*�b��I?6)]ln���92y4J,�ZE��-��Ʈu��iv��Qw�:��E���l���*�I\��TMηa�y���ĉ�����������k|��9��2��oP*?+�]ޞ��Ç8>w�di�+��7^����	��0�{��x񹗭!������EJ­��% �Nܙ�A�<�<R��Y޲2!��4ҡF�aӶ ��m�*&��詝8�c5�E �9�d0�&XV��g���plx�����C��0j�n�� �F� ���m�b}������m9����a�q)0}Q��a��	[.��r�*M�a���}s�߶�[V?L� f�G���9L�����~�>� �n�c}����]���Yԋi���n�@;��{S�\ ��������0��>��8+�j����/p|>�;.�t&��61�	^���r�;�X٧��=�P���2��u&�}Q˜8}m�>W�@a��F��W�T���;\M�hu����|�>�K�����y�����>ɿ�6L�F������-�I2U�n��C�O?�<6w�Ĳ4p�f��r�&0J���S,	���y�.���4�}��g˖%p������!������p��j3r��5j�� ڢ� �~.���K��8�\�e$����i�$:�@����\ F�jp��i{���9�S(�hd�jg� 	\)��S�m��$U`J`N�{"sV�L Oϭ��tG3�']S�L5y���wU�� �����,���{T���a�ޗe�5Σ�� ��Ԝq$k7<2��ֵTS�s+��+�ht:4�z��e�J|��}�']׶��9~��H2��6�w�\�Ͻ��6~��7^���_��|�S ����ұI*Ol�^��c�I\^^�s�OM�-[�0�RC��������-+җ��	[����5],�<4��:��2�˫K���PX/��'W�������������NW����K���O�ap`�P��E11�t��GD��	���o"���q��Q仉pl#� &fO���F8�e��L_x�={�9��Y�Bj�6�o>6x��E��t��������?������[���_��� ��o��%���:��Kv�N=⋡�-���޺��Ӄ�����/|�J�t��lr����xp.�������h%Σ�7�t�7o-��w���q��a�w "�*�Q���:�q�����)��N$�v�X���s�M��gｃO=��kȦ�(e	�����7��<|��g�a�v����x�<\�3��G9<0��L��`xh K���P�ڨ��scs�f'F��9��0����0�-�Ӟ�[>�|><\7
�>�����Ea��D�T5�*:�;w7Ш�nؗ`j0o�Ƹ�]|O�rw]Sԑ�T�s3�� M��\�}�r~\~v�Y��L.��	KM��"Q�a��R� �f��gN�gG��I����!�bu�F�E��ˤ;N7j"��6�[��� ��w�`���/9�� :�!λ��zba�Ut��E��4�qe胡l�yL`��K.Rx��N�aP�����y��*R~���=ڬB�6�/�o�ƽd��1��j��%9��\�%�^�5�j,o�b�������\��6��g	�����Ъ�Xjo�@�����]��M�������	+��z=&'(�٦��}���_������F<�N,�Z��S����C�$�ʕ�u�:������QP�Z�Բg�"�r�.�*���:����NU��P+����0	)L/������̈S�K�]��p�yP=� P��]�K��,2I�5J@7�V���H{�Q�H�C� NLҸt0q.�K�>��[7�p����.�{K5�l�p���&���-.bu�Y�f��186�l>c ��uwo�7���������P��q� C� �Ql�ְz��H��#�:ǼiYU��;���:K(��f��_��7���Jg�����I�BT8uk����	��>T�N�8��5�Sѹ2o�{�j�sm[>���VWX(��sY�I2t^�� � ������-NѶ�Y�p��)�F�n��H�ԅ-�f�L��2z:�����ͦ�鈧�'�:����t8u_j>P�QvS�����T�F'$���[:��:O�����c�2szOz_ί?�-\�s��wt=�BA���>Ai�d��`�t��r��B�wn����q�U�n�AF�\�^�Ȁ�g�����;��!L�*�����i`�ʇ�;����� �/�]c��[������>����2���o���_�Ct�7�3i��΢�P�1ȧ�uI��tn+��x��%�V��zۇ�K���9�w�,��ֿ�ܥ/!Ul!18f�j��ۈ���q��x����x�C�����#̜ǝ+�01}�z K�%�?��pd97w006B{Ѐ��@2��P"�߇��q���h�>���8{�"��Ѡ<\���+�F�[!�Ƌ_|���7xx�o16���c��P�/�����<D��25_؏-��)�t-c?26n�-��ꍏ��5|��b5��ǿ�����]�a��U*5����Q|��{�{�y�b���'�	Bv102B0����8�����d,�1�H&D�4��{;OF15~���a�J;���#82<���,���s�mlbfv��n�X���P?��!�(D����*�x���P��{�&��pl[5��VE��M�[����$!��;���q��9�+iM�}h���[�u�6ߋ���B�wP��s'�!�����A���!mY���ɗ�F$J@�Z��\�OA=4���{z*L]^��3�K��]�f�o:ƉD�$B���j�=tj$�����I	�`Ě�J��Mڌ��C|��/��k#�O��Y�pE����c^�L��Z��ٛ���%C|<��q;{;c�[�Zo�fb�s��O{v�s�s�H;�+|Ʀ��3a�&Ւm����/M`u'G�K��w���j8����
�� p��O�+�����~��˹>>���@�a1���ݮ7�$�<ց,�GLWU���rq�`�����M�R��!���t���?�D���d]�^Ru�:���㤱j�z^t���:��iZ�px��YIJ�K4L��Hۍ�T��F�pAf3�5����(�*�}��TB�;C`Ql�`�����{�hܫ������HC�ćWަ�o����� V7V�����M�@jF	EX��1�����A�"���P�ѫ��؊��������OR�Q���{��#�`��)��"��vy,�0��=c�>�:m�2YL��t�����ʦs���f�2��H�y�����<z�f?�QG��+�gm�����C�1�S���߸j�I��-k)lo�Z�GFSٲZ�aT4��) e��\!Wm�OMO���6��!���&�Lm=�3�!h�cӳ���wv��iXuF�j	��"
ǣ��P8n�Y3�j��d�|jZ_2�;e�T?��SOaei����0"47Op�w`NqlbKK+��������l�?��QxxW�<���!�<���.v7wq��i��;{��������޽���X{d��_��݋��~���8��б�>3��~�'�	�[%��@����[�;�2<�2���|���<-?�m�ĵ�w���m��������F��щL#�7���5���� 'Ng�n]�b	���~
��w���z�-^o@T.H�\��7-��η�����hg��`����(_���{Rs��Q�t1 m���,�9�t��"?����ߩp����-�J�&�@�֊�G�[��Fx������~|1��8���h�����;��PϷШxpƭsuzt�������k�x���XOm����t��׮X����1�c����~T��h<D��F�hK�x?>#�?Hm#�nc4��R/�M'����)چ:�C9��� ��g�/�����hR���\-��"̵�qW�����r�� ������e�����.�C�l�����s[ip->u�"��iC�����0B���B�*:�u�����s�@��8Oc>ڊ&���H��� �I�E��Q�@@�)zW�~�D��I��N��n���e�(^>��s����g����c�-h���t������{7_��cS�����w��w�rZ)Q��弩p�'P�:��?�2uZ�^-0'Ǳ$O�Z'���� N�?I{���MDg�H3�R5��r�o�"m��c�D��F�~�a��XP#f��d��eͤT��"��|I���0�q<V5y||��s��p8�*��.��l4gǊtuH�Aŷ-���͞V��L�Ѥ��H�#Np&g���L�X4���>��+V�� ���o�~��^�Dc�MEy=J�ڌ2�lTF�l_���=V"��[�?����Q8f����|�۷���v�xP��Pr\�#Y������b�pD��Z_���9=;���aw�FN<������,>��MTJ4z�v�V���Eg��J��"|�o���}��FϔJ�5���PcM�ϯ��\/Cu��I� ml�[�0J𸼸d�#�ge�����G����$��I�5��$�h��e���:04�����\E�|j��u���)�T,��k*�&um?>g���
_}�U�n>L��T&Kݛ�c�=��=�7������R�#bj}W���0UV�;��%��N�ww9�iUM���u��*V�N��ַ��+W���t�W�\����"�V���^�ޏ���ܼX��	�Sݞ]�?}
�C��E��|��ٶl���*A吽u����:�+K�t:]�z��A\���W�"��#�-����te�KwVz��K;�e��9@*���N	�L	���:�fR<��3��=ol��ν���;���^����Cցo j%���#I�\}��?���=ˤ�	L�������N���ԉq���G��S/���.���L0�?0����M��%��FǦpb��]:���k(n�����Z�3u������}���xL�TD��o��l�#3��;~���]F&GQjv��vCct��~&�|n7oU	8�m�_�<�kWoZ6>���p3��u�O*\�u���I$�_A��b��� ���v��SR�~��"� �e�žcs�9"F$����|�>����1>���7#_�t!���ɱ���h��@��tʍ���G��Jɂ�b����F��C�c���I��8-Hld��/-4��; ����e����R<zk�*��#jT���bKڒ~?b�����X�AIOF�T�X.Z@x��$�Vis�������4�yt���?�O�����
ܴ�a�C��\X~��+���~��A�ͱ����h2a�v�;�hgv1C;1"0j��Egv��R�y�ӈ"�]4��x�S
��fO�C� �/���o8 ���歉�떌]�X�S�����6I(�甎|���@*?7�c��]�Ϝ�=?��T��Ћ��<�"�V�1Dp62�o; Fz/>mc�*x��mv��e�&J/}�JFԘ"�$N�:�ٹSX�-�A��|wg����S\˛�v�*#��=���׍�U�#�*/q��6e�fӶ���_����w�p=>���|�4�o���\�p��]ӛ��Ѷ`�F4Kc�"2?\QF������FC�b�o3��<���ɧn�X�R-g��C�t�8����MP��
�]<�2Amg��wZ�5mE�F��i�<e�}.�ĳ��Õ����7�i�I���㧑<9����m��	�g���������<�}�*����ݤCG���Ν��ϵ�G� ���m`m��Z}�4��,�YP��ؚ[Dk��Kp�o8��V����Nҁ����	,T�gʪy�f��بu%����O� ��r�l��J(�4�[�H�N��R'�逺?m:�ϔiT�O�'�"����K�O���ehe��Y�����_e�^x�|���vNGmZ�{gs� ��,��&݃�S�y�7��v�c�мj9��G��j��-i�"ʀ}�w޶��Ň���s�{���Y�}#�@��~T�=l�n���Kc�p��8�J�޹oY�8Ͽ�����=2�~:9fQ��'�M�ĉc������,\�L]�N�3Ϟ����P���$�@M�O��u'��#� �sf���ÿ�3�����O���,�`_�����׀��#1/��ʓx��ܻ�.>x�oq�������Ux�f�2�x���U>�L�"��ۚKp��6��i���X�����5�e��� �N��.^}�/�φG���������_{���eȬ<�����%��^�8&�Q&���%ȹ_�����q��o�0N��
�n��@�`xo�.��X����R�x�?���ql��p,��OY�+Ujټ���!���L����['s�:�}�!��F9?R�"H���-�;��'�!�h��G�l��v�v6�'��Vl�?����
�Z	o��Ѽuc�u�.ئ�V	_?�!~��C�]�X����m��sIҐ��"��P"���x"M�(�g:�k��P�P���a��>��5�h��A�t�CN��Md����À�P�#B�1N���Q��w�`\K
�@kWD���F矺�u_a��j��2ׄ���k�Iq49��n��7�^�:�<|���TRElo��8����q�+��q*0�%i�bnl���7�n����繖 !��gOю�Yp�M0�.�Z�J�O��D�m��BZ���4����{��]�R��W��ϚȤ׬�e�2I����7D�Ġ&�d�I�����@����a��szJ���Ό�U�f���A@*I�J�j �mК��k[��&�S�etN��\]Y�����y�ߥG��B���Jvʼ^�a��|�����V�n����萑���Y�.=acP��̾��/@�c������|�¾x��y��.����<Q�a1u�vC�"���8�*
���b~�
i"��A$��F�c���1��U͸�~���NT2���~#���|e~N���渐Ul-�aƀ@3H ҧ�XM��)��A����~��`�69A@���M�a�O<�ݭ[pS8;����w���(#]Jᰒ���&��� )���Og+��҂F��,�����*����2��To��4��݈� �'��[YF�:�?����5���tG#4t��>2�p�<���p�H]O`MY,�ިg>�߫Z[ؓuK� ����Ԙ! ��u7+C(�% ��A[}�H[Y�x饗��2�����@�:w�{�9S��9�e���9�'�gH5�����=��F}��랏:��y΋�/a��=3)����6v����8��K4��2������!������M��s����w蔕����SzTès�'��)�1�8�r��>�f�'.?�7^{��4�sd�9�Լu)��9�s�9o�l��s;x���/����n���"wQ]Bt\#�̤��X,l��Q?{��Ezws'�4�Y�:�䀎�o���f���GWo`h�<����Oo#�Max��9�6Χ�Eˤ�����G�p�6�Wpz�,J��� ��A��A)}����c#�w��E".���`���ՃH�^��.+��76P����:�ν�z��w4�ݻ�r3 ��hљ�x�Ln���j�"��ڸ��g�lF,�
`s�8d������_�m���q���?�;ps��6�������6�.�3SQ#���X}��w��i�*���c�����o��X���G�/��>g�B]e�>��;���ne9��$F����;�W"��b렀K�~�3{x�����I#W�K�6�^DM6ѥ��.�D N����񣪣+30��B6�Bjk�c�6Xyps3.LO�3��mRx(�ĉ㧰p"�9�	>{����\G�l���B^D�)΋�5��i��������;(���p��f�/҆�2���I$�t�lTf��pw���1��B��ˏ �jg��3����ԥohڎ@�ն�iѽ@�����z�j�����6ZkZ��i1����>:AWOw����А�?��J�����d�r�%�%�kq�a�vӶ�E5�������и��w�^���W�de4�<��I?�lv�V'�9�F[184��?e�\��B�k����oA���C�����kд�}����u*�j����1��d��pv�f����:>(�x���5F"�F��+m�>ۼ䠊�)�'hNS�n�F��i�1d��>l��[6Q��Ϩj�"Rv�	��d"j|�j��1�-��mld���3�k�������P��*��b�$\��í�[�E��]��N��!R}cc��:���,:<���(��}��,+٥s�x�F����8(`��1l��Y��@�ȷ��-�Ռ�3y���ٓ���:X�����e�ҩ4B���A.��;���5�C����=��h1F@��:,x�hW[�F�УGQ�Ϛkx��Z��qԨ�s	��Q�W�O�9�#���G?+�{C�C�K�R�N��nbm�
���Q�b��?y�3�@�M���b���>�O�&��9쩜Hj[Yu��T�Ԉ�i\�L!`'pۣ���H���#��j�J����}ƶ�u�;".�,�t :�5յ��[u�tTI�W�_��Y�9{�����Q����x���`_?
�i�;]�-��셳�������m,Ju�o��XVtff̮+ \��[.BGX�񜞘µ���S'qjv�����z]��v��"ܩ�_ϡ�"�*��߁?��V1�7�beq���ך%8]ܽ�k�p�u4:-D�=���.��^��Yjarx������� Wi ���o]�zLL��|p���Jt�-�3�V�4�?���0F�e\7���ku|Ei[�QH���(t�۵��/<�q��ĵ�N�����p��XY��h�֪��,v �J�K@��E�u�&-��q����	:Y��m�+�����h��nj���B� ����x��,��5LL^& �"A��E��=v�M�M������0ױ[�{X�X��Ǳ������ϐ��̹������fD�����H��0��$c5�l��x��X��a����8�t]���"�:��	v}ѝ2��i#�}�g����S��c�{�
�7��1���._�X$��`}���8�O	�%����ORU��=�?�7���1�E<��!��~	7�~h�8��(��
v���i�G������W���x�[����Qm�w(j�Ej'�`�Q
��0Vc����ڗ�	�N��;���9,���}����"�0������7aФ��v�'��n�X)|w$�c�j8Tm��:ǲ���b|u�ʖ��҆&���!Urц�!E[$��J�c���P��yc���!h��)r>��lE�.�9�Ã�Ո�1�M��F�˧��X���TY����LMG��+�ice���ḱ]�Mee��U�-su��.Z2�Rb���h�<��%���F�&&q�v�U��x�����'sp9&��jŬT:J����A�&�{�rɄ���(�u{�ET���2�R�$��H��N?�f���M0C5�A��
�O����b0���}���]��e+� h���V-�t��(�k,�C��~m���|Hm�ȳ����\z��Ew��<�+F�.,.���8�..��Ed�B�~:c~n4�������au)E0ڴϿw����K_��޸����|�/�����u+*,f|��e%�"`�����c�|��wDD��#��j���H�9|�(�%��JQ�h�R�Ae���� ZM4.&���y4�G�4G���)�&@�L�@�>{�3�5eu^5�h]���^`P`S�BG������3�۔?x�[�P��^:z��Y=�}��O�MEY�'�x¾�����ߺǣ�e���Q�U��m|e&u��4���L���5���n�]5H��3�y�1�����ᦥ_N7�����L-���5�8��pОI�6�iiVgs��o�S)�~5�}C�q�j�
\����vo���e��c~����'{n�	v�W�"P�Ԛ�*3�e�F�z!��d$g�f�A��~�+`�W���L
���k����Y�j-Ē#\�js2�s����W���q�)x�����|�te'O��\�v����~�����?{��k�)Rc`xtش�w��:�S�����G�c'U�����f��"Ю��#�J��A��*O�T�V�*#�`��m�1����\�|gd�d�
U�?�όc}m�@܋��1,..�܅��" Vk}t�m���w4�?L�炗�Lo�p-082j���->�]�N�"��|���Z#���p
�Ç��+[�s������}a%�$
]	 X����8A��U������J�t�%������;F�U'�QP�C;&��?GYۨ.����$A��}���w9΍*�F�8{b��0Q��`~��+j�b����Kܼ�6��Wn~��@�
�୥u��c}�����6mI�_�S<��p̻�9>�_z�+�^_����8��Bfg�׋�g�-"��r�xV�Rx�ٗ������.�+��=K�9r�GP(�TG��1���m[)�֨�iz�[=.��g��>#;f�H��13��OvD%F�R�Q-��~8�# y�6f��Xgr�>ln�Ac����g4��[G���ڨuS F;|�uײ �oh�b�s����Yv���qw��79G�Cݛ�}^���,�ѵ�r��+��'��n��Q�y�F/F���>\�N;7n�-s���N'�O�����������<����j�{��M�S�F��7	T:&�78��)�b��سHndp�X� &bġ���b,�J�٦��f�I�Qk5~�*�I�794f79�LD��n� �ۇE8�L�
C:SuP*�68:a]|-~��,a((��yu����u��K_Ư�����N���+����E��ǵ����9	�'F��tlf�WM!�Hz㠂��1�^|t}ǲ����1<2p�w�����/��<�ß�G�;���!>[�R�z%��V`F�����n�m�Q�WgwԢ\i�Jjjue��E 9?���˂	4���N���E㱵�c��2.�@
��M��m@R\�22��D���"}Ӫ�A�����>�!��w7�v�0�8	ܨaH@M ��ߙ��@�T~��ǖ�3`�{[���l�\`V:b�:�U#��hS�:�@#@���u�1�A�
lZ�_<n�ӵuϺߞ�MO-Dϭ:H99�e^��h]�;�|Ţ���'�mcm���`��xl�=�5�ۻ����4n��VFU��3�>������Ҷu��N3�������:߱�hU��{�2g�� �vö�	'���~'b~��&
�"�}㘽�
�!���Ǩ����{�&�M��W0��"9�H�i���{�N�Q�H�؆��U�����ə�|�}��# �5�㪫�Sp�$�����[�����E��]�y��^:�Օ�0��keq��6Hg�`�����u|��5�uL�ޥG��v���M�:��[A2��#}]>�`܏Z9g��+�Ǫ�w���TsO7O׋p D@�56��Vى"�gb0F����,�,��K`�� ��G&����X���������ͱ��`3UE��B ���� �-'R��"H�;8E*�N��%P����e��zW$�F�	�������M\��"�7�-p��M��ͤ����C��^�?`��S�2��Q�m���)���C��>�
���xp�ML�yi3CH2��%�H��C����
�1�G��J1�K/�҅)\��U���@��v�RBH�R������F9�b��WS��cr�<
|'���� ����8���@~^�U���G�8wl�m�����1����eL�]@ؓ�S�Vκ��}b�u�����y�O�����Խ+�����+���bv���h��A�v>Dպ�M�9�]�}C��M͕��X�+Hg�P�083�Z�Mf�P0�_���$8g�-�;`r�v6�vM�IV9^�EQ����닫�Vo0@N����kX�Q._ОM�m�;�}w���Vс����],�%{f5����5%�B�ےڃ��{��������/r|>�B��5{l�����ZÁ����������<N�nc?����H$d��;[t�4��}�F�����h?#�7� �X�G��Q;8�Ւ��`��)q�5DX�EW+g12ҏ��ti(D��n�>:���>��@ۅpЃ W�^����<.�;�H���'!X�|S�P�n��1����`&U��{Μ�0�s_� �N��*�;��F�~��\۰-����Y�Վ=$�m�9F�.�Ǜo�au!ɾ66VL�^�G(��!u0��x�s����˗���۷�zEF!���L�J��8�}J�4(��	|鐁R�J�L����\��֔��qUVM`I�6ێ�Y�:ʰ�oe�������e��#�e�G�r�:�"�.?a M[������H�w�nO�F�Q�- �m_5�h���:,��i����ʎ���Т+��,��!���\���({D�-�d�)ꍕ�ODq|�������a��!,�fy���	|k�Jc#�b�9e :���/�;�W��48>��%N8��o�k]�ʆ�Ξ���|�����ǡq��`����E2��T'�:������g�?0���C}Lq���]��!�>�J�YCy7�ύӣc�-���-�x���z�?��Y?>��DB���,�=�;�(N>}h���S������<����	�{��宮oc��6��6׌�(x){-ՠFӅ
�$!=���0�7�����{'ꚗ~�<:�f�B� AC�B�>��rtT����Z���;��Cu�:	�ʈ�c���hT��`��1<Z����U���O6W�(���KOb4I��L!�9��������G���"(J����Ipf
x��s�|�v7G'����p29h��K���e'��u0�@�Q�IL�_��}��;���;�W7L�S<�Eڶ��92 �VC�j��d�ָ�Z%{(a7����s�X�����
����{��w~g�h�����/�;x� e�[D� h�t��8sb�������	����"N�ϘԚJD���`0�s���~̠��6���M���f&1:��� ����%�~`'NL�之�����x�q�9uwr��֭�F�d���ZIq6J�MN���&>��+�/e+��O�A�����#u�� ������ KeM�*�=La ,��R�i3K�b�xm+�1a��)�^�|Z�jt�IQ�[��P�5�pyͶ�c�N��S����0�!ы�S�%� �m��]�y�ڨۮ�>k& �m��ΐ2�?��i'�k]�w�+��S�<>~���u7JNNj��NO=�UF�ø}cw�.X-�3�^D�Q_��1Lb}u��#�fYrL4�*�uy$��T�:�>3N:������px�f4YG�Q�+��~U'*�=�g����� ��l}sW���^�`�F`l,�V��.��d����)����T���f�b)�sT���@�1����� ������b��ᩔ���/������C�%�բq���C��s��-���δ�zlz��ǿ����Ox�
söUﶵ��QF���R�x�s�Ȩ�M���m!�	)&�;�<Am�m��<y�l�����=@��Ω����@��������gM)2�������b���d("��w�o/��QVQ �|��,a�-�r&j.(�<D& �Mq\3i�"	���v����"r����=Y������k�)wn�Vn��n�����2�+���ݱ�n��lqnf	���j8�޴#頓�Z������>��b'�~� fg7���A䷳�ѩ�&c}u��j~��ػ[z��X���/��?��Ձ�q�\�d!H���k���|��/���P�n#�b"�1uq�}@�k�h��8��AL#h�[81<���&#t�6x}����U��W�G��
���K��t �����ݭ����� �5��k�Z�ߥ&8�O=�2���E��� sh����&�����R.t�����Ū���u��D>�?��{�g`�L��w�m�!�ݓ_�~iB�̉kt�]S�hUJ���g�,}N^���3�񜺜~C��s�>+��z�d��\�rَ��!�D�A~w��ކӃ���]���9���x�jn��vܦ1���-w�-d�� ���F�l?9C��b�o�8W=����\>���_D�͹Xh!�`繗����~�c<�{�mJڙ��~U;��Hխi]K�W5fU�E=�����y�����8�k���H���1:����y �D��ܦ�\����S�V��Յ*����-�:9>MP��I��'�#��	�{��aff�� mA�:����<z�x�N;�=9i_��
R�=�V�G�SW������<���*�<:~��z��äs5��/���IN�����m�]�x��p6]�V��*D �iY�;��x��m���$��5��p$i�rg?���:Y��!�(6����}dino� ��SP
�P.�s6UM}3���.�ؠ��3`�zm���S�{�C�5� �����B������j�:V�u���o��g� d����	>�E���X�j&��F������s��I�;EּH��.q�'q���	��!_�±��C�o#�4�閪%����+��y�4��̮<I2-?xhQR6�4Ap?k��C��-Qu�T�t<q�[uۚV�0xa��R�".^�G��=��ٓG�wo��҆	��34H�[8H-Yנ��%K�{zp��)V�Wq����Uݦ�s�3���Tł�hӠ4jU<��%�y�?��_��y1>9eJ%�� ���/>��;wq��A�	�jgt�z�2o�X�JٚK�g�~� �b?e��{6���տ�F�G>��� ���Q�N�Ki���������2gOڶ��mӉ�H����j�Y�/G��gG��C#t��,jKU�L@T?�Ϗt����V�6�^�"ZS��x�r9���[�P�U���TM�����uN�H=��V-���mS���D�=����������L�S�}�+p�˖��VΪ�"er����w��CAٺ�o~�7���w����O�����'�۷���Oby}���ը����8L��ݟ���!�� �h���.�R"�eRD��n5�[۠!|bp�)�9�&"Q�)v�t#����Zv��l�T�Fyo��p��˱���t�p�H��	Z6��r}�0A'�4`����X�n���؎�/��b|j��q
�����>�Ӝf�Y�<|����X�/}�cߏ�G?W�AZɡh��XYĘ�i%	2y�BN�Zk�T�%.�"���m�>LJ�6��f�(�v��12!z�}��a����c�Ѻ��8����o�p�*��\k�h��h��8~��Y˞�S/eAOy������eS]�.:����� ��v�n�:xO��^$P����a�Գ;ε��u�z,��đg𼻓��\�z���70<2I��Ɲ�5S����,s=�@"}���3���)�d饗112�H`�`��Z�h��\:�b��L���5��� @-`x�ku��/趚Ƨ�?c6�ν<��'�	�̱��n� ��`-�@C]�\������͟t�� �юŇhUSp+hBTkh*�~��SHM N�*YpX]��퇫��qWFL��-[��V��7WB$�k�Ӝ�L���RGV���\pXW�l�4h�<!�y��²�-���Q�8��"�r�mL �sE�k�Ғ���0(LѦ�	8��"@+�� E���E����&�|�bM\�N�$>��z�J�ڜC�]�75̨�0���AcR`@���X<B!��RU�����ց�ǔ4���}|>��z�Q*U�1i��FO��L�࣫q��,��(�������k5<N�
n��Mk�w8��n��x15uF׻{k469Fn	.ښuC*�Rf%���P��L��b(�,�"9�V�e_Y����i�hM�KUĜ��T��`�<��(T��I��1��)��� ^��}��9�W��}8�nlK�VQ|�������!�ǧ�I��p� #i�p���u����׌cp0��Do���E}��;�m5B7�ݦ��Zݖ(t(|t�XI������E+͆��,�UѴ@��i��*�slzƶ��I��phkS�Q���pɸ��1��4�S� MFT ��ϋU5Q��j9����MDc��K_�L��s�C�=u�@��l�>1{��w��,��l��w��zJ
"o6m[D[��G]��$JO[���� ��b�=�`ᾁH�
�	��!��l�Pϫw�h��� �
�E���e�Sf��ݻV�#��`�Ϡ��|�hYK��^|[cE��H��]�VjvP������t�������.�ލ�x�W񕯼�M���ݏm�Ru�� 	�Jrog'guK[;����N�9�}�L��}KίI9t��y����&��u֫�,����1h*�ꐺe�-��r�]�uW���F����,[Xd���4M>KF�uMP:C�~��jt����Z*����]��\�cmI*��˯���$nݺ���3%�F��=��w���;v3�|^Vn��A�?�D���kG,�	u�j���^󘲳��!���[���Y��&�s��TC���E>>=�����	�p�憽�d"n $���Gｋ��p�6kv�$��~�}�N�ǣ�[p�~������=+U��q\+q��m|�)[�����
�j��=20�50���]�I����_\����o���� �c�'P������[w>�]7�4���a��<��}�yb�e��ֶL{]ud�?��t^��nY��,]����=��a>��"��6R;71u���a��
�NعΞ*�!�>>���A���Z��p��<m(;ڵd4bAp�k7���i�u���������5�UjM5�T�j�K���j��i �I����q�=f:5y��M���r�ֱ�ի�S坤�m�H�2��~�R����d�JF��Z���t[Y Q]�.�sM�?%�0F�U>�ﬡ@���L��CpZ��[8@T��^��BƂ�w:w������!J������xD�q��=IS��\:�
�_�T�y-1_����f�VO�X]��:�` .�E���(�
��� I���`n�nX(� ?�����������F����%G^�b>	�<�T�2
E{^� ��&�6M[X�k+�897�Hԇ�w�`g}� ��Ss�8%x"�(-"��I�ڡ�*�U��˰��^�A�4k��}����b����0�n՟dѥ��<],4�j��!�_� 6fĠ5w%��7�TO�̃xa��d�jmF��"����bss�`7�}���Vi�O_��%��>� }��n�@�����^}�-�;������k����ee`�d@@82�O��k$A����	�z��Q�Pݸ]n3�Cʢ��A%6��	���;u���q�g�L��գu��m4c�k����(���?���)#�s�����2}j�еu��IRj�/}O�����	��zGu�����ʦ*����~��T�D���?�X��k����s��w݂um�L�X�=*����A)���,Ѡ9Gr����&Ev��=;�3�<�����¹�g��k��G?���������j F�"5���~�?{�G�o^�|�:-<\����	�:��vt��]��
oׇ��@�<�!��u+��R���l
�y�S3���?��ܽ�:Z�� ���)��˚�a��M7��;�S	�Z_:ƛ����F'��p�{�XY�M�k��[[����ڇo��H)_�lw�����>�Gc�x�+�Z���w�`z| �L��C���N �lh�J��`���!]��\�.^�͜H ��%��1#�L~�M��W��Ocxb��e�ʵ2�j�IrL�Hs�S��ɡ�nb;�7n�瞽�6������/|i��׉h?���+0������-�akӓ1��W���D���~�'���8��],�*	B0w�8�zk��8��E_T����!�������L�1 ܲ����X`b�*��>=�,�8Ϡ*A@q���v!���{|�Yڐ,ǈ`�Y��y'�����Nr�0��T]z@>�
��r�U�y���8�y]%2]�3��d(]�����5�����C@`�����t"�u�s�dK�R����r�A%(�6�ۺ��V*�L�h�z����	�#ШT���T�P��
����d��ZYU�a�^y�Q���Τ�jYnTis��{MT��y�,ej�AR�G���$";*}s�Z��}D�(Қ͖���P��d5S\ǲŪ����nr��3 �h-���Q�s��ɓ'8a\���Z�l�>�dJZ�j�k-o��..a
�ԍ/�f��u�<���Ǐ�_��\��ϙHĽkk���%l�,Ӱ�Ƿ�ѯ�?e���G��wsQ�at�*%>6�Ħ�	��;���p��ϭ>���m����3�-��V׹ ���a�qA���sED��M0�NG�Q���e�$k�#���7�۾h��c�=�-���us�/�й{fzL0�� I�hY�(���h��.�h��V�X�\�Ქ2e�$J)��
$"r0�<�=3��u�~9��n��k}�i釪�����{�����ח�j�V�v��Mo��1#�n�k��x��~��q97�*7�:w�p*�6A�d�|�FU�����SWqb�$���4��hf��^��8�g�}��k���䋸��{XX��������������W~���{��^�54C�t���е�	8��(9n)fѦ��V3�E��1�� �իW-"@u�`"P�������1)���J��ڶ�[=���z�iC��
E>{�3R��s�ԝ���b�LR-����5�.}�*B�W�K���L��w{g�@�����zf�>mD�4���c����T�O�'�o�_`X��zM�,0k��;m��nnٽ)=&�g�KI̩XI@B�Q�Ϻ�+u��V�m�S���AUr�~�x�����'���?��~�0s�4>x�->��X�tfr
��o~�@o*=`�7o���/<���|���� D�u�	����&���;@�s(��V<lGѓpC
K1���M�č?&�^W����|������9���9���A�Ry��W��lcR�O��ѱ!r}��VJe�t��t4�9#|_Ƥ?���x��ɱ�9j�+�Ъ�164���w-5G$�xσ��a��o��E�`���6,�tbf
ɸ6��O�5E��j���ϻ�^��Xd�<���x���W��|��?crd���5Wv����Q,7����f�+G.V�֬��}O|�"�XZ~Ʉ�|��`���D��4uz�Kwq�����E�a�d�G��E��up(��o_���<甈���'�gp���s�6F��JyQȊ[*�5:�t�Di��>o��.�߮�ُ|Sw
���9T���Pz�^oغW֣�?j�l�����o���8ù�������������֮a4V��6�Y�R�c㏘��E��h��jU+��4������%둛`-�GS%��_N7�R�NzY@��o��U�^�����������jWL�O��$>�o��&�Y�aK1��CC��TQ��e7�]�!|����?��Z��Y��uD�/��n�s_j�����<�wz����CD�:��+�����w��
���8���M��v���c��z�f�T�󫜤����"����ҡ�G�Dc)����=$�X�j��N?J�����3���0wj���O����9/О�`O��]�:���ǢY�H�[��ǭ��Ti�a����'9֋u_ �k=*Z�� Y0"�����)%���i
��v�"pPb/�����7���`l�4�4��+�r�N*�NZ�W��~hulW�i(��bn�й|�6A�H[+��x�0���~�	�+�׵b^�-X�7�$c�Fp�ڈw !w�"G��eK�6%� �Z�b�b�ˍ����,`fz{��u�y"���O}��.N��Q��A�^v�����~���_��������5�����Y��:�D# P�R�Ʀ�٨������'-�:7��i��ҡs��P2x���f�VN�_�MT4M@F^��^z�ޣH�q|�|v~�W7EՔj��%3�bރ"���L� %�f�nr�`ߢz�,Jj����Ң�U5Ǽ��[&����!p����y���D����[�" �Cc$��8���=��Ng�Ӊ���A_��CFP޲��f���;(�3C4��o����CS˸p�~�o�m��3��\�j2z���籺��_��_���E��-=fE9����x�������b�T����:�����qc�নNz�j�Y�&T3mm͇��!;�e��t8�Z��=�u%��	h<���Gx��Ǔ��3?�%[��jN" &3�F5k��'O�`s��������ܶ5}��_��h��?�y0=1�9��6���q��02<esHuT��$�v��~��
���V�c���@:�n8��n��\*�n#�0�>7�g?�>��/r�Wr�6��s�?C0;C篍�j�6����R���q���K*B�������E��!#��S�)Ԛ=�is:��JK��&V����g��_�*^~�u��#$28u�,�x�6j�?�����E�����/��E0��>�����`O�"Ƈ3td�Ж���<8��(�B��s�����[7	�È�&��c�������5��KB����4��V�`�h�߽���,���Ϯ����`o��!B�i��<AR��?��P
�\��yM,@aĖ����F�YD�F �)[�I88l4)�~�X)`ݿ�G�`����{�.K��igE5�/����+@���Qk��h�M�C������P�;^�'�����E�b�N���Ã��Z����L
s�'y�&�G-d�|F���p*�'�f�HE:Qq���V��$�\��`��("J[��{�n��.�c�x9��}v������(qZ��"��Dڢ�zVj�R�H85�6(�Gƹ>g9�!,����_�p��;fsU������i��<��$H\5IX�"�/�$��_MY�߇"!��<��?��@��Ҫ��P���*-F�t.�^&8:e��R���alt�ˋ��Xr:�M�R�o��ŧ>�94*�\�!��X��w��@O�@ܰ���`ay�EǇ|1�1.�d�O�sd\|��R��K��J'�j\Q��7�Y�E}��nT�Ǔ�ˍ��3�[yǢ!Qʡ�)`om�~�kx��s��q��C����A��G��J)�g�y�sn,�[��5��4A�o���l�X��7���m�7�7�[����/���"}�;��[o����	z�U�2˅<����J]��j�>6E�=p��SO�G�>*5KX}�"54��nf�-�uW
%� �}��X�uN+��?�Ճ��R^98�C:�2𠴬����t�ի� ���̴m���.�;ŔŋF�Vc' '�x��e�;�>�����!�:��I3ҏ�*GTE�J跻�+:y"u���s]'�OX��"��G}�����*A��6�쮷��u��ovO|��[R��������3�ŋܞ�`z�@����jـ�׿�u\���Eb�6�0;;Oÿ��>fQ���}`�Q��<�����k��K0��9&)$}|݃&�v�S7wq�s8�H"� ]_�׫�"!.��35Z=�m�c7�9�_�j!9�E�K������u̝���t�	Ӷ��Y�ޛJ�X򻼆�-���/}�`����rK�Ɖӏ7�뗱�~��Ғ��Y竗`���q�EB�їE�Pd�n�9sGH7��#{F�[(l��]�c�(���v�6������� 7¡T�6�ӧ>����u)�k_]�uu�w�x�Oc��5�=+�Kg�>V�z}��W,-{ga� `�s"Яc��0�W��@0�@��%@��kϿ�<��
���3�8>��O���5��!�/�M[V��O�ӟ{��ȋ�|/��{�ċ�F��n�M�թur�h;2��o�EP�-�UKX�����I��diC�� ȸ�tךQ���%��XZ��;�{����-TGP��!qf���jBW�	�9��/�q~jsggqm�}>�=�+���E�szq���|�"?j�n}�ݱ�*u2+����CҮC�"n��n���Rj�eu}JK���M{�
',�ע��E8[ChW�,�4j�J�k�Hs.�k��m�C�d%�I��Al�n� ���	t��!I#��`��Jm�^������h�:�Fj��(�.d5%�n$���9��mj�k�1�P�J2�h��]����I�Mg�Iۨ1�e�2Q:�,'����I���8�ixCi\y{���):Oy��� �u�˵�LGY��\�����ė�3x��/�O��a}m���2�>K����6�� <��:�"��V�Q��P��Vn��(
�*:.�X��D��l�F-N����`sg��7�S\\~$S�zК�n!32�ŵed|��XŚue��5��4m�0��#���:-#�kSW݊���(����m��ǹCQ�/�En����K�#�Ս�/L�n��7���	���[z��&�4�J�D���p,�M�����n�8B��5����A4ª��w�6��i��Y����� ~��[�p�"b����o������O
�?��Ϳ���]Ckk+49�ON`hp�" }e/=��Ĥ�B!3D�a�ԉ�6�U��D|������me��N��4���ȹc�#Ic�����D���q���j�h]x�Rz�j�HJ��h4���#cc4\i����ҭ�u\�r�"v����U�"x��<"*������S��}��E���i�kvM�I��ʾkL�TE���Lr1_pRՊ��j�)��p�Ϣ�|��~���_�x�����II3r��j>y�4{�<���ϝ?㤳7v	�n�}��3[�ScT�����K��ŗ>������6�	g	V�^�mJ#!>,r	��'�m�5��� Wj� ��F2��(�7[E��q��m
yx�~�T�ԊHg�wm�VA~��A�� ��Af:�F1���W���xp34e�q�ҫh�U�T���a�����kH�b��F�1�Mb�`�Q�����):tc$�5΃�iH���Na}� �H�󷄅�M�!�SB�`h�����L��|�\�Cn�A#�Ҟ�*El�T:A�oc��͉s�XYH9�B�P�{�����>�����^y�u��a|����y�sOr���YTUv!@`��E1>v��.j���k�x��7T�oj>� v���n-ܱ9"ȯ��������s����������;�hur���K� ����6���˨�����811�ՃMT	�#S�N/��(~��L�E�1E�Z�a�BPڳy�y�QT����+�I'k�$���I7�kx$�ã-:���-?�QL�a��aR	��^�����H��#S��������[�����cm��B1���t{��ݎ5��KR�0��5x�>�w�Y1��^����4^>W�q�:B�k��U�31��k��t\�J��h���@�5�t5M���ȳ/L��똛�A1_@�Z��X�@^���������/:��^G�:�E?Eg��9'M�f�a\���������S�UL�KY���*��V��1	���+�9�X�r�v�]x�Y��pr�4�i\Y�>����~H�)B��=m#����X]��Ż���x��˸�9�̳E.����\��������B����xx<��@�P�#J��5�*=�:J��?q��Pg�*Vi:�l�خ��O�0[��&S��瞁�]�����1��y0�jh�[L��X�[�~(�@�SǙ�	���o("SAh�����}pQ՚��(�E���ID������������xznJ�yh@�"SH��X�r�R��4FEb���7���]�d&96=DO?�O$��5�0|��6�<A�4w�gf�a�c�Ԝu#�w0JK4�b$������*����?�_�[����C��y���op̎��%�����)���^����E�@���6�� q|�՚���F�!@wLJ��Z� 
Mn�;���s��Ua��V�*���������	�כ֌�C�����>E ���R��J��)�c�� ����µk���+���M�-b�'j�\���JyK5�n�[�͌�"�|֖B�8�w]�7Oİ��F �"N����98�70�x���"�Q�evf
�Iq���OP)��9�vu#���3Y�k���w�kJ���]����{`�{p �[�n`����?�E�$.�Y��А/-܃���#O=�k�ns
�ܙ���2�
.<:�$�Q�kM��CQ�U�[sMu�>k�(s�D�\w=���q�(���182�6�uST6��ܝ ����-��F/�X2���e9�ܔ�M��\K~�����g�F�;�;��'Q��$ ٳT`(Cg��s�M�]�MN����{XF4@4@���"�*Бk�v,u{g�:2S'q�T���1�|&a�K���	���"6rU\�����]��FKIl-�����%4]i\�q�k�>�ɏd����C\~�Μ��=�'�����?�4޻|	5���p�N����ҡ:�A��
E��:7]�[4�����'XR�П�鷸�����B�����_�7�����71j����6�Ƨjk�u�.���{�p�qE��;=���u���o���J�^O:ۥ�=�*&�N�njP->���3E����ɧ>ʹ�"hX�Hz���^cA�'�@�jY����Y޳;�.u�Ff�-���R���Bt$��$����"a\[�ґ�t����Jâe=�4w�Ƴ(����ϝ���z-
(NL�z�e)�6ר��ֵ�m��A�  ��x(Չ/ۡH~,����[�&-�{-���S�9N�fv��}�/����\煸�N�*+�H�g@�Ү0�!{W�Y���������k�c����v��^ٰ8�o��Ňb]���t�j=/�3��ܸ�x�c��+?�6N�=��'͌��'����j�=�8�����בH%1�y������mb�6-c,��tT#)%�`���=��yx<��@����p_s��X�%��J��ѽU�K������k��Gx�$�\0����H��$��{�a���P��1o)֭�Μ�GNݟ��+�41n��F�AmW��H�q��(zM�쵝�J��'P:*�&��6od�H@�Ko���-n(��(����F�].��	�;N1=����߼E��C��zL�&Ë��J�7���Q\-�����%�z�W	pR���s(��ڹk]���%�v�n������M���[Vsv��y|�q���8���el��A��!���2�v? ��:,�R1�堁/�&�gu�;���Ӹ\f��+%;��Ș��Օ�F�351���e��)�"�s��ju�\z
���7����8.Int�����$vJ�������Tt�͚:C��S\ngO��QO��LMY4U�.��p$�A�q~�Xs��-x���o�R�֝'����[��j^�j�j3P#��F�"�!Vt0 �Ef5J�*�o��ƶ��h^���{���4	��|�;8U��xw������}���1���\"���^i��J��P�p��[�J��P��O}��lC�!L�&���|�~�J	��������4�]���)*K�h��'N� =4i�D �:z1;��4�	y�&�_��1�>*��^x�E�[���wW��،M�IG-�������ͭ�sD���V�?���y/c(��,�2�s|JR� ������c	���[�w�
N�࿒��@���� \�\��Q#��F� /���:�u��_�^~�?�8��
�=���~�����;5����<�(ԭy��:d��on,bz�<�G&��07{�� �{�.�:Ry�:�Ϟ���_�����T.�k_�~��~��p�`��q��9�kR�C"5'E�Io�*=��]ϥǰ���
�2��o��7��?�%�e*�=�s��K� �Ȑ{�/�"L�Ԣ}��]G�����
Ξ�#�o�C��S�!]�x)5?w�txs�"�?�Z�O鐠�e����l��u�4�Ͳ�,�d���(�#+g{��r�-����`��B�2禫�3�';"�ߎKTIF+m5x�Jr��Kn��:�]�*'�ص�qe����Ɂ�I������h�)e͵*.C����]�+�k$w,���K��BDصHeϹeNIu�]©����-j)yGݴ^9����� ��r��;`�kKk��k&gNѡkc��`eu� 2�y�m��?�忁@�$6�KX��bh�������sO?����6^}�]|᳟����:㙌]��4�N��ｗ{H^��x������^�������~���&�ALX�f�AV� �K8#s	���Q/TФQ��,bg�6h�&�G"3��&`����F	4�ֱ&gM��x�o܇��u�9��eעY��i��E8<�sa��Np�5��P�a���'P8����Or��E�����(b(����q��=�Ν~�+w�_;B*�%@I�MTrr�v�	��ȣǞHu�3�󧱲��kWp��Y�C�s&���z��������?����ϟ���9# ��c���K(Kn����w` D֩�0�潛槩ƻ�ާZ�ݧc�SS�q��j��[�~h%���%|���g,o���`���R���1w{B�G�[�I LTgi�;75�8��I3������U{��@5��@�Ҽ�p���z�6�J͹���y�]�\;�W0���r.H_�od�*LWDr|lҨd���mdJ�;�1+-�S(����(�Ь��C`'�o�r�O�a����8��P����9DK��|�����sv��<zO?�~��7o��3�@O��r�F���b��A�����@2����(�W70?;���UL�z��/��������pX]���fFCV�.5F��>�swj8�9�'��G�8�Za����F���OYz��%�Қ
��{7�N'd6�(��Z�y�C��Z�ǲ��r3�#15��\�s��r�@YR���ZMf�m�F��"M�qbf=u�r�5���Zm\8u��7w�	*��yT�#X�A�3:/.k6�L�`t(Ҥ�RB5g�n��d��%�'@�sS���5Q�����$ןd������!�:n-~����}��QO�²5AK�f�\�~ź`���Ӹq�&���b�v�������p
��}C��x�G�b��"�t�O=����8�z�����������hhW�^v�b����:jy�u�g�(j{�P���c�b����1��E���6�x��7Z�BO>�(A�4��m￻�����Xs]u��R�/p_�Y�GX6U�}~���~�^��������l�C&��T`��wB��{֏�������8�ԩ��U9��?J;��C���iݩ�����79F�r��o��=T��q���ڏ�-`�Zt�c�]	�+�� I�l�G簟�q-v{-,�ˠ��be`*���w���	����ǆp��*�� ~�����nUP;�`l`
��'�B��,F������A8�zd5f�������ߏ�S��F���rʇ���?�x P�C�R����ɕ	��g�q���HMO�N!� 8�e��/��W��ܞz�W�Ae�.�<��R7���%��L�I�U������o�Fc��x��:ࣿ٨qA9�wF[ �M�oۑ�g(� Em��pJu��!R�8q���{���K?�ٙg����5~���t�mn*A�V��BO�8M �:��F�#HE���E4>dj 1��;�����ow0j��k�n�f#�v��	��EnGF!�ֻW��/�/<����(��?�O�A�1o�h��9}��m��׏��q�*�	�D�K���!RtF���_�w�pc��!3�0n
2�J�H.��뼟�m4������o��R$���VoZ]��1!����y]+s�@k��~�p���\�r��W].#��kU]����m�p��t�S3%E�����Q��u>GԸ�����i��9�>�:�qݗ��Z?d]��%v�fH�|�MD�0�ܡm4"���T/) '�}S|d���Hi��/y6ۈ����&y�y��������%�Ν���X�cB�~tr�PS#cX]�g�d"�>*����Q����$7NE@��Rs��l[�O�����C����-����*5���q�Z(e��n��%|�<[����6���?@<�܉|�ϿAp[��}�A��Oq����>�RAܻ{ɺ��KC��3-��:��=�9���[��2���
ؼ���o�i�#>:x�N͔1�\�A�P��i��D��v��&7?~s'��A��63��B�k��@��_��EcT��T��eS:�|�<���[���b��_�s'���[tz�ߝã�Qw�m�O�x�T� ��NC�y!��
����W�6�q���{+��UR|^{�q�:ma�j)5������r|���� οx
M��ڟ�����^��˭Hg��v��T?�/(e��g\6�bvP���n���5�Vn HX�uhrs�� PDz5`�E�T�)����\[ZG*9��ׁӑ�ql���D`�>1r�ӏ����� ���D	�N�O��.]��U��h��Yǀ�qD��i9���sLe���v�=�]��"y�unǽ���4m����H=�*t��S�q�����qD��|��^�tp��g���z����"nq�8u�tv���U鴨��O�G���o��=���/��8ܮp��օ��"����$j:Zn)��#�8�H?��?c6u�0�f�X����sn�?���C���
;G�K	��	L����bzv���.�e�]q���y�q����Π�|kYd�ƍ�Ѭ��	;���R�zG�r�Np��5[4�.'B葞e��S*=g�[�=�D��j��E������N�I⭷�X�X�@zw�LU�j�����R'gưAP29Ӟ(n�ZĔ5}�x�W14L@xP@"4�C0H`�^��sS�3����92�/>��ｃ��{x�OZ=����*N�9�m�o�����W����_�����������w096�?���⺣Ǩ�h�%��IB@�cݵ2�2�2���畢k����� ʀ�L�#lשMT QT<Q���o�0_X���d��QjVR�"@g5DP*��n�An�2�����h�|��Z�ǒwJK�.�m�ޣH���U;���ר6�{��4��X�׊ 4ZM�����uEu�\�:��h0x?e���L��Q��|��}�;?�zAEMw	|Z�N��pp��)�,����}{v�T���:�L�G����O�n�o��������	�:��5>�9���+cwu�)!Dx�9����0�E�S��Ωx6�T�Ƒ� 30�@<�͡n�LJ��QT+M�U�fW�p�Y�����~䏲��~������q���x�(�A������V7�����s/����㘺+����x�	T	��<ב���D�:��T���z$QV�����b�8<�4y��>�܄>��s��"�h��"FFƑ�pm�wjXީ��g�@�8�{�`i�[M%�00E(P�Gn��033�k�6���\?������6yM!��R��ܪ�q���L�ǉ�8����E�t�k�~X�����������7߰����͍�i�lW���Nm��_x��|��1���=�q�7p��(�����d����;���3Ͼ�����7	�8����U�N�	��:wYm�r�.���>��^���<85_(I�-�G=���S\���86�ᨐE2��O!��(t��$���:?�95p�����5�i�:l��q��n�y���{N����.t��np�	�~���y�9���~Nt��f�I�Zm�����W%Q�T N��"d*+��^s2>��C��;�������Zj�c��ܠ���'j�Ï�l�[�1����-j����"�Q:H�T��V(�{�w	��أ�08:�����@���}nK{���X^߰��z9K��4����eL���XYG���:�}��t=���r������く��kL��.�'��XF(~�gF*>J�����Qx]|�O�B���*F	��n�D+�kD�͈Ȁ���&Y*VMҭIw �3ߐ����ļ�5���z��F�M�j�����:@#PV��!��(���]�ȏ����7��WяJQ�]�^�����0�N��Ϝ�a�Ʒ�^��h ��n΀k1��*R�}sźD=�LM͘���2�GR�ٟ�<�\}#�\�p�`�n�4q��� ~�w�^{�G�ş�2~�W�;�/��ի�Ym�U���E�K4��B��,���#N�M�v��լ��8�!0�����6�xy��Ǣ~�f�X��~��HO�;NT���-�'o��C��`�k�~:���6�vw�+�xL��k��Z� K~x�j a�嗬�D�W��pk��6��e?��:Dܪ�a�W�����om����@�xաs	D��,%'�������&f��\����%E%
%�k���ŭ�Y�;���Y�=�:����o����|�*������u>��%��	��(T��M�{y�7��Y����A3��*�\-���ԝ�M6���g�F�����aQ�ݷ|]������D�@-���V}V��-L��u�`zЋo}��&�+��(T����x��k�]b�kF�<6�@���@�����k �ɹfRc=�^��0N��ȳ zM��t^T�)Z5��:��=nf����P��=|�A�D�\;Bם���D2�6�<�7����r�eT�6Q��9�BK���|�6w�|��N��3�X�avf���������-ae�
v��hc�19���&�Rv��H���i�b	���e�MAC S��>�J�3�<���#�!H{tW.�������uxuJϞz��{���D�k���S�.b���ѧ^"�>���BV'���M:�x��kʺ`3����K�143�&�|�pdN���e�Γ��1�����e�r�dk%�)g:�YdQ��� '�gi���+��@���D�@�Q���%��_�_��ۉ�u��ܯM�O���N���#�5|Í�T�bM#��9u:�֥�л��rS@q��g�g���{��qٍm)��V�u�rE��
�K���c�'�]�2&�v�N���S�l�J�'GmM^������k�`�����P���/q��<�(�G��F�Ο�6eGt�P#U���kƉ�����'&��bn[Kq:A=��V���ٿ���C�M w�'��%p�J&������}�����J�`ݩ7n-���)n6>KC0\�r�'?�FI�@���֚���﹁��5t\���ۮ��)#\@\�h��-K�&��Z��S��7:��_�Iqu,�k5��h���Z��r �=�)|�����#�6�Z�����a|��/��)�&�o"��_�a������E�A1�0P1A ���W�Jc�o/d�ZjB���4��"�L�t���@�#Trj�p7?X�?����c�����ayq�I����D� Q�-���X�a��(0P���J�j�9�>���� �����N�kQVB��<A�@c���ך{=��guz�4HNzPD˝f �B�^H���of�(k3R]�@� ���_̕,:�)uL��p��N0m�:�`�"��u2�X� �J��dT�W͐q2�~�='2j�
�(8�1g�"�F@K�4��z-l6*�$m������ܑC�����w2�J�i\��*z���,��^����p��K��2=;fe�r���b�6?=�N��d"��ׯ���Gqsy��U�?A���������d]:Otum��|ar�	�TW�1M�R�
�H��(U\Ģa��R��������u#��R���ٓ�qs��`gN^@�pu��'��i�. ,�gΣ�?B�`M�Tp�a�}��ߨK�P��q盨SQRtS����t�!NC�q��}0��F��s�M6I[�pQ�?�Q��[�آ�$�}u,>dQ�u���
'ǧ��A:�{� �	T�x.���}�Д
�H�߼�#������4���8�����m��v[�w(o��dzĸ���O��P�Z�b��(��]}��LG�[!��4��?�%d���n��W��X���@��dƆ������� r=�yN���=$ l�y�qzt3�I#�\h ��U�(���~$�n�⦶$�8�d��u���˓k0��� @��wXĬ�D���~&��q�m�h���h2�����Iw���.��u���>��bt�W��&��um�N>�t��S�h6N$R"=�s� �J�%g	4V:�ߚ����~M�@�S'�O!�x��{rY��q4�}�,�y���>��C�h���.J�N���v*��u�R1TZQ,��#��s13Gۿ��xb��L���ci��m�Si>�����O�K�Z��(�\kB}��/�}��&�[퇝����x`�¢sn��/�I������+�&���49)wh��Ѱ���|��>;q
����1�`f�G;���L��j��Уb�^����M�dڥ�@��L4�k���*��Z�ύתg|~.��X�)1ʹA���`d^��'Щ$�,�ЭK�̃P0j�s�}'�`F��(9<��A7���]��B9����~�6*ɐ͎�beu׼V�&QK/_�t	��r5��2��͈��p}eMz���W	��_}�����:�$`����,��E~K��FU]�2�}�#/W��Ƭ�WQ�qJYMj�(�K���hp$�BIS�8,/�մ��+�OF�m�6��e�"�
>N��<��S�6�����l�F���j} k.Q͍>'C���EN�&��i5��B{�#�
��7�H�5�NZ$X܎:��4�Ƶx��m3�S�36R|1���w�~5�E~����j"-R���� �E�{|E�����^�E�4�/��r��ϏY�ЩR'm���������!f&',�M8���MW��������΍�	�*#�z����������+�$�)?�I��u&Zi|W�&p�t9aBn�~I�W9����>���ַ�[���m�{�ߪ�! Y�/⚼}�.��C�x�8T���������p�5b��%�Ii۪�6c8Q��TC���"N��j�M�P�=��J����m�-i��5���aS7i6EJ_��]��Y�0�ǳ����� ��m.���4��5����b�YC�ǖ�1?~�����b���;����"��5)�"���[�`�'�i˼(�
�]��R��� �z>gc��?���h�$��k"���f��'~s�3���a�Ex�+��*��=�.����2�2	�Y$J���^֖a��*����]ۺ���íf��I{	.�t.��w'�,i��.a��H<a�Lƅ�Ҹӆv�c?�B�W�pk:����ϱ���>���hbkD�H��=�;���.=�28~��âm�ij�����sá�����K�8��� �}�TmϜ�)W�g��R�}�N�qr��NT�w�|�=��}(�g���q-��k`��=W��
E��k���6�]�,8l6��J}���z�!^�Y�!��#�?@81H�\�qh�FKѫݠs��?����B����8���]���;��pv[y�]S��Gk��E����Op<(�z=���5�*i�ed0��_�&�^�8�Cܘ�c����҃)`��M����{���>�9,�z�y.�@�L9)�p1�CI�m܅+�Db$f�u���FΩq�ޤx���y�]o�~3�ۺq;F+��P��j����$��uU"�$���}�jۢK��k�Xڔ�ڹ���t� `Ǹ�>�%.޴��������(D���pf~K�ܘ]�ΪQ�鹋g�(�0�)lT�D�!LL�Z�8�Fƍ�nqe�ӧ0ɟ��e�~�:�|�*��L�x��sH'���lCJ9*�P���#�VG��Gq|~S2�O��t!wi�&��X�/^O�m]�n�Շ)�,�1��ڲ��p�$�$
ư��o���XZZ1���АLK�J� o8�n�ao��jLr�yK�e(5l����(�Wu���	q�ϗ�Ymq��,T�(7�v�M)�XZѹG� Uz���G�V���@��C����mrj�����\>k�ǀ?d �
��[�YH����n_K�Cc]��ٙӳV���N�ɄqPf��V��5Ք
���a�ܼS�X�b��9E���Z��3I,�/��_ `;@%$>2~��{cg�1=u� 4�����q�|��uY78F]�H�]q�scW�8�9�J�i��3粈a�S��%����t2ε\�p��x{�σNA�iғ�pۤ�D�n�p���󂄞n��+��9k~7鄎%��1�qx ]�����TG�\Hjmk;�{��؉7�
;C�B�(���(�rk7���"W!7Ab�����Y���;=��;|�'�
�tk�C��w97��;O ��3��S���7>�aD����o"�#=�#�}ۛ9ڼ�m�r(.�{Ě�Fg�=���K��(ayy�F���E�ǦO�O~�:�!>/�@��m�k�n����vǍ��k4W�.��G)�1
���j�Q*�E��&i"nq�&�ʪeX�4�͢�%�t8E�NgQܔ��ǹ��!�V��)M������r*='�*������=��r� ��0w����r�b�@���
T/���N��*J}A�:Ի톑C�"��Z�Ǉ{N�r?b�S��j�{})Ϯ�*k�2�.�ٮ߈r ���_+5�'�I���Dur2���Ub���J�G�9�ة��EDU�Ӫi�m��dƪrbW���^ۤ}��!L.��b���f������Dq��c:z;�[r�r�D�6���ݢ���A�:��U:T�C�Ȗ��C�Cl�����	���u�W�f��x<M��Í����˘�*bt�<Jܬ3Cq.��'�z^U������0��6NA��q�/��Z�f姱���w�E�^q8�E#U�D�RS��j���X}CP����o�9)z���2�n��P�dh��GW���A2,5.�F����w��1{5ܹy��(����x]]���G�85�!H����y�@���I������3�hCE�4�411f@���$	����i+�(�����*2�|���)�8||j9f�8n�0:�n�{��`5�q+RP�5�)ZɃ�8�-&��hZ�ݺu�v��V�j�1�a��d��	�z��7-U*V��] ָ���	|	�����ad|�\zGBY��4UI��U��G�AF����R��k������b�h���c�L���"W���AQMmB�
F����'XS��6�ѡ�9P��ʤ,$c_�|-U��6E�8uℍ�����(�V׹��G9������ʅ}�,�2o�r�|�KL�p�m��O��[7.�X*��9D�=ޫ��>G�13y���W�b{�]4��HĂhֺ��}Ku��o��[���趚}
�K;4@Q_��9\��H������3�T��R��/&�Ӽ^��U	�獺(�OP��XT��nc�B=�26}i:�J����8��H��<��v�9!�Q0�-0��M�i Q��6��q>�B�=nm\�w$,EwX8Dx @��`����g�r۳H�ɑ�����:@$�0"�hb� j�sr �PjM	�6��%��������f褵,8����"@K+Hg$A y�eI��
��.�;�H�6D<��h#3t:����\|VGhw�=$��p^��!��3������p.��y��Z�s�BӺ�+U�`g(�8�t�Ă������a����;Q��ׂx}5��M��S������M�N���\�\Z�"qx;_�
��=�(�[�5��+����-���Ee"܎�RtVK�6k&2�R�j����"ܵn����}����Q� �:�1��JE)궚b�}�Au?���t��~�Pu�:��zv�� �c �ObYܤ�/)���%��9���5��k�8l���W��?n��<��_����R�BS��t�W��#9d"c�U����mB�)�� �S���i����:CC��)Z�C�7s����#{V��0}���Ɏ#�n�]���dG"V�#���~�W8�9I�� �����ӳ3!kB���]�b�_h� h�F�����ϕU�@ �4W�q����@�{���]���>�+���)���v�ƨa���@1��υ��L䧞���㶁Տ��7H�R<��#�?~w��\��١ 
�������SX�ZF�+c  �^���%��c\����k;�M��)#���Scp�\��,��rc95n�Z��Ƭ�N�%OM=b��(d"Q�A�A�ó�p��n@����咧ۢ!Sǟ�8ӱ����qC�[�(�����&��A=�07� �h mS���a�R�����Ȥ�P}��70�����'	�&�8M�o�
���oTvz��c)��*oXQ�G����-=8D��v<���}�� ���XM���>�1��� ���E�t(��HF��I����u��&�u�:�25�Ȩ�}n���DQ���M��R�Q��'�B.�7��zHטh����4�jEL;�z)���i���Y�� �J2�@R#�!o�B��`��'������:oI�����g�V���q$"}�Xܗ����"v�o�W�E��B<���o�[_���٫7+�T�$@,�-PP9*r���ԓ�p>g����g_���2"C���q]�ư��a%"��il�x��F��N�(q}��+�g ]��P�6`�qG�Z�R��P-3�q�(��r����$'�9�#��ӡq���=׉�PN|�W��4n�
��*J� �r���b���б�@%qx���@1���a� g4>f(S�aL�p�]�l�e\��p��W1�F�����s~'�'�,�`�C�����Tllٺ������4vp�V0�R=l�/i7΁XЋdRZ�txZU�d1���$O5�9�t6��[d�v��{td���MT�?������C�N�u!W[Ro���G9�z��5&���K��gu��A��CU����v5�>���K�^s��]�(�V�c�R5�|�>�I��VB|���ju9O9�U)O��wr8)�n�0�tJ����0mE8	$;&��5gJ �2"RE�S�X�J���ix�سi�~KvOB5��K�d�ҰR7��*5+������b�_?Rh�:n�&���Ng�ew���po�k!c٢����(�f�ʮ���&��h��� lu��r��|h@�x��?���qC��?�:�G�8�����騨L�mlE,���������FI���(���{[N�I&��9��;[�}�5���a$S�Z_����� ���S�CVܭ�񼵺��U4�y�^�Rai� FR=T�a�Wj�8��袘�]��D�+�s?_C��&*$�t!���cg��~$�+FO��!x���:�p!��$@#�TK�#1x.8�,o���5N����g�Z�h���;j˺�V���6���\/�����r���L#ki[��T�֍���e�Č�9DS�=y���ʢ�
��䀆����㪤ºfA�6:�	�z,jר���ПN�e�qp�!�j��Ǥ�k��N� S�F�QA{� �i�1��)j��PiJ�҉Ʉ𡋏�����?��x����}�:��,J��>�J�y�&�^�s��ܐ^4|���߭bf8	p�"�jܐ�k��G5w���kK�	̟�&D��r�$�y��ݶ��n��X
��h:�y�O[Ί��"(�K�Z�4i�TPT��F��&��t!
Dz�nR�T���Z��C�(�@P��qO[]�av1E}�,�*�VAy�s8�2�ñt�����^���S�_�=��6�H���A�`G;+��K����n�������tu;}2^����JI����)����	 ��wYy�Xz�Ͼbـ:�_�C)9T�����%q��N���V�oeZ�%ڳc']w"�����U�z&�~
Ѣ�=5ɸ�Z�Ū��6�CKH�NCe!U�Ey�u"��N�c��"�Χm�a�H�8BǃS��
;�*7�X��\��W[#8��V��1�5sM�����+��?�5xD`��#'�U�87�
���<��A>W�����[k�-�Z�a(�/ⶒ�|���\�jF��	޸������m�âT\{�P���6�k&D'�-�G�[� ��k>�U9����E��7;U�t-T+��1�ւ��<y�~-aNp�m�[[���V6ѳ&�H�c F>��8���� �����+�Գ@����k����-uˆ�s?�����R���u{����
qG�l��[�%*�*m�oʔDh�6�R���Q��~L[���Bs�!�J����5�S+����I��c{0);b�T��9^J��ukb�G(��jE-��#'��d��0�ʱx��i:�-k:�X��ə�)ls����>���2�	����x����~��:��`cs�'Ҵ�u[CN��kܼ}zŇ��く����$ܒi�f��P��M8}t� ����{[8��f��
:� 7�H؀]��Bn�QWW�!`��d�Qi]�|�4��>���@t~.��h��6}M�7�r����r�&�)�I�*�C��Uu8>W$�a�J�)��3�gj)*��Vs���Lu���l��C#�Ƞ�N�)h����RݭfeQ���b7V:*����]�)�N�V���ԙk�-.�v׀Ti�nѪWz$u��C4���EezNs�G ��C)W��U#ؠ����Ep*�$/X�¹|�<~I�5��>�Dۚ-$��+UfZ�j��,�qr��*��c|����/b����?������I�mn�!�Hڸu��2G��ߑ�OQ�tY)VuI��mo�����QzY���">��XZ����+N^,��#���&�\ko��k��>v���6+4�:��VX�/$����z�N���,vJ{���"8O�R��J�����40��5O�.m�Қ��m�R��xo-8Su��Z����U��I&"8�-|�R�ẇ��y>{�Q#x�U���z�:�:�a�Y5�j�S�<��`Q�VǢ��|�H������j3�b�pô_���Q4y9�(�ܱ�MSQxS����]�YAA����`���gC�f��	���^����y�u[D���~I��z����V�F�q�>��Z̙R��r�A5s��.`��V�L /g�cum�r�&c���%�u�=kf+fř:b`�KС�]����`g_Y�0�s��9�!C#��H�;��`*J�X=,���k��̼*Z���
�'����f ��(�a�c����È='=� �AJ���|�/�2�H�>��p�b �����W�U���3#�6�֠��}T�R.v,Bۮs�B���zwש�`j�>J����G��q�׎�j
	�|.�}ŏc�;�X�n?�j�rT�I��ఊ"�\ob��..��Ʀj��@��j����y	�*y��m6�����"�����~{�TF��v�H��Z��B�u#;�i&��]��ʟ[w� K 90hMgj8�p�L�ʺ�]fC̑�9P��^b��J��7Q�[*����z���)r�8�MIr�ҕT143���_�����0���s���P �bz�$�[������-:�v�q��M:(�\r��7����s�8<�����x`P�B]IAő��#Ҡ6�I�%H����A�R|G{��`����K�YI����F����P���n����T(���4T�j;�P4d���4ƴ)@b�[�7����w7��S�B'���|�5�IE+IQAu���A*_�i+���ڴ�)�nI��Xe~���&Z%�Rؾ_c):W�8AS:����ޗ�Jv\��p��T��d��Tb�hu7��6 ���7���Ѱ����/��7� ��[�5r,q(V��M9�!���NDf>R�v��� �W�e��{��=�s���4�1���w��Z�l;6�-R9�x����W򐮮֔��Q��S�l'����;��sX��$��	�����g������2��ܗ�ѕ�)(4+�E�i�J6l����]d:;.��<�nXQ]�h�~#�o�!�
�=?GZee6�O�Y^�N�*��nP�- |V��Ԗ)ìh�JN� .�{zT�#p|~"�����k��gZ-��}h��O��?�g�5?���ʼ����G��=S�FjT��F�s�W)ej�m�v2X�͘:J�=��]��`a�z��!��4ח������'��~h(�*��-ֹo��es���߶W�jNeN��W������~M�����'�}��W̳�O̕�~"o\^=#_��ș�S�`�H� �R5��͐Q��=�V���a�7�b,ٺ�����
���XL�_�慢"?8\�����-?Ŭ1�e��N�#P���}IN�C�ޥ��("�1�[�6�v� ��sG@08.ȁ2��F ��g��g�+6itB�����IM'G|���&����[�lq�S:=�j.�?0��\[�v�����eaY�r6�������W���s��W��������¼t>#_�]-Y8������ �F��0TL����2Z��e�[r��Z �9���W�N� :��*� EH���_rM�2�'/��}���������]����Zr����@�Q�ڪ�K$�B9�p�|l�|zHa=�[��<���{���IQ_�"�z�=x�elCz�/~�6Sį=x�\�,̇������e�e}���� ��\�]����1�@l�E����lx�Ĩ��<���"�Ӏ49����(*�gXlk�U��^��<�|�f��5z|���fa"� �)�Y��I�?m���2KO��#��믿`>��Z��er�af�������.������dV��̯�g}��?�o�_{@*ͯ�c��)�zm����О�Sv6����b����۪��=6��;gfu�CJ�.�M�9=AO�h��|*r��xqu)�n�4�|�ŀ�d�Űv��!}�b4K٨'h�$�wA5Ӟ����}#��!��t���k�ݿ�
L1�T��-�(���|�O�^���n��F�+��+�����mP���	6N��+k.�IZ��t�
�vq�5�!a�	bh�b���ܗM�-s�ʦ����ڎ�sr	`&�kUpC�<R ��L�T;�7#'k�L�s6�F���
���4����	���X��@te���,)�jvBP���c� M�n��L�	��#�V�w"A�`l�7L�@"��ť�����������o�O���ݻ�)��g��`�C�ظ���{�H|������ &}�k�<�xj������P��P���E:�|"��*"R�U	����N�h �h8������pߑҺ-��̻O��̦	�|� �w2���ҧ8tK � ����'����Y_�Nݘ�Ֆ}f_����[ZF�N���pr�r�p"����D�(Ԙ8�A�$��d�����6n��n�[���%�{�F���d���y��������a��dCaۭ�S�����T �%
��V��DC���5*z޳ՙ���q�i� B�D�9(��鮬}�jM���h�BBX�:��w�����l�r %
k��Ll�(����jYdp}��6>�Q̖iM�5*�Q�����M�Z����>@��y�K/�X��������gzs��b%w�N��F��r��ȑ7WW�7�N��+���ن��=Yw2G�*��Rb����)�3�o+���S������L�V�R ��ښ�9:gfX�w��_�&W��/}�X,��� ���b-@u���R�!�
�D�a#�Q����߈6�R{��|6ha+e[x��QY���)�?��N ������'?��y�ч��k�ɱ�))<�g�M��V	��)i�@L߰Q	=*��8�'L�#S2�Q֍��A9���R�TR"iW���'���B+k~i���TJ��o�&�����%�v�S^1�.R
�9X��n���hu-�]�n���a*�Q׸���{�y���*�������3�/��>������ߙ������\/�K擧����G���3���;�<*�����tb~�:�B�q|����խ���٩<1K1�Pd+I���W�n�=��}X7�ě~f��O͝��V���YI��
`*���Ǔ��N�va���U��,)x|�o�d�\�Ll|�D�3����J�%�V��e����Q� ��1S 0	����TaM*�6�6����T�(a׃�I��D���O.\�1���׍��� ����
F-���Z�Y%*��b6c%�U�Gݹs�Mu:��KG��T�r�d
�<�H���1$PV�^]�LM��-��я3�\��{�FS�,��RJϨ���gYՌ&�(�����AL(D�ߋ�����nn�-d�Ҟ��Ĝ�&v��6��`L0Y�"f�յ��`��X.ds��7z|4gEv#�w�ŗ�o����G[��7���'� �u���!".6(D�Ph�B��<7��	%4ZD��+v����A�YvZA�2D	Q!����� ���Sv����l��I#�v!�Й���#8�����	P��;�
��|��'t2��~l�Njs$뽒s�#5�{��-�4��NAW  E��)��bH˼�SH���~(�ͮ`q
6{D��9�xc���m�:�P��Ne�f� D��P]]/x| a"iT/$�JC=J�q$�Y"�F9v5�,�I�ߥ�0ht��>���f��RK�J�-[!���nɹ��
n#πn������$Y��`�ڰxL�a�B�Nu�
d�	�Z�fFO�2����} �o}������	G��3F��g��4ʚ���s1m��yڑ�<��O/�QR	2W����x
�S5��X���*�+XRqaH���T.
��0=;95�W���/�g�+s�؋�ʼz�E�A��Sa���\O�]���&�W����5D�O�sSώ�6r�S�A0}j��<=�R���_m��N�J��|����ʓO�������+ڮ���6t�VIJ�pm�>p�s<XFx�ݽcNOU�԰W����B�lPΪc�G���
B`�R�\	~�Ɯ���=��C�{F�J�ж�7*��QR<[>�zaHQ¨{ �Ǟ$�n7�
O�Z�eO p_-/h�`�_{�y띏�~�}�k_3/���=����جڅ�Kc�<}W��4�����U��g惇�b� ��8���(�$q8���f����@�X�n�MQ�I=gA[�-�e�>~*�м����o��S��5�DJ'�tZ�c��BODV�-AZ�u(v�T��,H?``�:���vQ�Ok]O鹯��V ��/�"�C~[O������,p���F�(��u�KeS�e��S^ښ2�QH�����JU����	H8ifbX����ݣ�U�m��8�a���q���,'���ߜr� ��H��ܜ�'4��\W'��X6�׿�*%T�E���ߨ����j(ǁJd�2xU��jմ��L����u�` )7`�
���텹wZ� �ŕ�G_�*�v����BQO�RhU��j%|l�|�,ssM�±����\
Py��Լ�f�l����z4���$=y�I�kAHOCY �>�H�m0��@�G�4J�$|H>/4���]�#h�Q$DT�lq�t�a�s*N	:�`����V�]#`��є��Z���bk�_>a$�{#Tn�ݝ�gZ���{
��D6��x��vW@&�T��ڞ˳�J��vZ���e84ʁ�%�A64�s
`��R�3��4�Mס]t�,�
	oH�r|��ǐ��*�k9���L�Ş�ޚ�O��:r]ʞt	4&a;0b#GT]c�_�?c0lӸ��hf��h	XɆݯo��*��&����_��fv�`A�U�c)3̈́��Яz��g��Ĝ?��m"?~(N��g#�3E�?h%�BYK��X��(vK��X* �9�rqi�X���O���<��j���e��v�3b���ʏ�Z�2�<�2��<�/!�9�K�hyF���1�Z��@ �7�O��b{@����N����S����'o9���H4�+HI0�mT�3,���Go�?��ӽv����wN�'�>�V�b7�s|�2��\lc�ك��T���D� {��9ҋb��Eq�8��k�-=ѯ�Y�`Tx�{xq�)1�s��o�n>��c�8�=p������8F�\:n`��My��8p��se��6�.�t�,P؄h�v)��¼��s�ʋ�8�?5�<~��#Y�+�K�y@��UqD������~�w�Z�6��템ѴR;�Z�r�H�8��x>�jy*jy�'��+��=� �,hA^�0U�(�t�?:X�� y��	�SD�*M�#X��	��B�2Jվgڠ�v]Erw/@�P5P�.�#��M�r!�{1R:��nJZ�ƍ�:��w��{��,�@.��:���D�J��P�,sp,�7Ү��V[I�H�ӂD~=n�	�b8��ia������f0Ǡ�Y`$ibh�1b�&`���"�U!�}R��+	0����*d�t�&��&�Λ��i�H�!ӭY�ݠ��c����@�!*������f��*������X��T�l�^�yT,�`���s1i<�>6�0x"�����'^(�A�p!Z�c�ԕ ����1u��4�FD�쩬�<8�X��TP�kEHG+rmU�l!�m��F���YCXCQ�ҙ�c������������J�y��U*Oqh7:D?�-,@*��zu�x���L���)���C<� ~��2&��#�̭
������|���MZ�nWi�'��{����f5�����͋J�`�����_Pm����o]�OF����A#Pc��IT6<o���uH_�TxD%���,y�Ri�s�
F#�2�� ^��g���5*�Og���8) ]:O��F�}0����x����!������t�|���|l��\�G��� #���x��/��(�����)j���h���!��"� �?��k�+�!�6s�F�Q���$�5F�B�Ey�˞|�Z���R����&t ~�y�}��DM� ��FNE�1�����ڂ�F
� x�vJ����?��hv���"G���{��{tf�Ip��B��b�h�AC-Иϋ�èRJ��4�|ÚЃ�-��H�C��ļÍY\��l�g���ܼ��C��Μ�~�������T����ӧk�����%`�	Eo��*U#�ؿx���8��x.P�oW����.�����]"��.j��������P�=7��X��Y��K��ABa����Ei?9�ɂ�5ɖ��2Uc����3�ab-4�q���*s��S^S�@I�L5FR��2�B\ޔ�nS2&��4�L�*~��(5tG�)��{H�Z)���5���ڰQ��7��e1T��7K0�T�j�1����X�	n�]�H�B���c1���C�O_I��D$k�:��f���y�?Zr�)j��GaId������t2qr/g�jyc��.{���=�\�+h�Ϯ�T������FD7�0�����m`��  �IDATk[�=yW���DY[t�)	b�F�E��h�D1|E6C�)����_A��fQ��.~/*Oc�*cp�b�8�?�U,�:���4
���(�!���ECh�59���>"�+��漢3�on�8�k
��:�skS����T�	�]��tH����`���}�m.@��еH���씧�?*,��mJ�9̲��[ߛ)uBL�@Z��K�Vb��Ԍ$��l�t��k��. �E�l`3���o�9��=PN�ݨ�v3 t���  P5�V��^-���A� /Q���>&+�q~��g��;�$�\�4�z���I�#�A[��߹������#�`)��xn�sf�R���\U��x݈ :��Y�I�4-����Tt�0׈xS_��� ]Er`��<yO8�`u��Ѩ�4�a��5���iBo�I_���Bj6**���֨z��A!@3��}ۍa�O|Ff�:�P����щ1�N'mAܟ�}�b��5�ɧ���s����=��q5�L��%;�T����c�Bʪ`mq\�M��2�9X#rJ%mzF�ص��8�b;N�LT�a{Iٞ���o?x˜�=�Q����`NO�Cؐ�>���Ē@\���8��x.PX�n�c^H��)��Xؔ��R�������B����daz,XR3��+R<Я�2ȃ�F5fPpA�6Mpc�On��$x��4� &�jsi�J���ޒ�m���~tI�ꮻ�u��p�N7Zx�T�wj���+p�q�Jb�]"�8t�Dd[�!0�Zyi83��e���5���w�c��Tc����oM3�%X�f���hQ�)F�
�Q��r/���) n;��]��X,.�3*'��{����O-7���j-��eղ-|փF}��bH�;mx-Dr4irqN�����5��^6��scfG����;�.J.�V���t0�:%���F#����N�"l�آ�N�l������i��lt-�*m8��j��K����	��W������F4O�.�h����h�ؒw�o�H6�Z*�nCT�*�9��������3=m�p�wj�ӳ�iX�I�a�zq�R�@9���e5�j�n���+�O�Z#g
�(����*{���ۙ
d�7�����y��[�� � ͍�`3hW���]��J�kh&A$�wVS�F�_���0�DiDҢ�(}���8=�X/����h�@.E�1���t(���|�B�dWR͏8�-mA>�!����$���̀[�<����ϥЧ�e�Js��n�[ΘG���Tӑ��@����'�ǿӡ�`M����_eA��{�y�m�}oU~�i�v-ǯ�nJV��5�ׅɐ=r���y�.F��� ��J�>3au����7tP5%\�Z���i�F�� �2��Uc�s�cSp���e�B����5-i(��~�vX1�ϩv�W,փ9:��c�Fg�s��N�|���sB���B��ۘ�e����)4�$
����VU���N���)b ��wCk�����^g��
���G��ީ�k�S�ېY���Y%��p���FԬ���f�Q���|,w�sy�$�C^�}f���C緋���	$m��,�W���@���$�0�FZ�R&t�M"�	��,y�c�Mf�ߕx\��e�X���T�|ĵ�3�%�`R[=m*��<���%0ػ����z}~��F�kN��u�h'�|Ô�aƪA�<w�ܔ&�ET��1�Wϖ���^C;(hUkg)=vĖw�~ Ռ�~���P����=ݥ�#E�О���C�[����sE �������R'�Fz��Mc�kE�2������4�C�f�!��*`{�4?*�����vmAr���aS�5�T��N��d{��e����|Ҳ�ɑ�G��u���(��>w���=�E4�{�#��b�um�>��@�ۥ��U �a���
a=���]�L�����	$Bf|=l��b��!��Z��w���D2��һt!�g�גAX�^��Ec?yjr�*
������!�c�y��Z��e{���p.Q��ooҽ���-(��g��1=W��t�y��w�.��¨����0��L��G��㮸w_�mS�F��)-*����-����=�{��nv6��j�4:�ȴ�������X���|F�S��ݲK���V�Z�ّm�I��~�1K�I�(�����:1y���q#�i���Au��D�I^A3O�U�ZZ�D�!a�C �_����>���.�ub����'���G�1��=�g7e-��
�8�c<_����ւ'­�ز8E#H�x���=HĔ�ꓱ�J�۔
�@-s��2K����^�RFy�P{=�d,����\�q"���K}<)Ƭ@,$����썙�9�E
wa2� aWۤ����B�2�VY-�iȒ|3B>�ceÆ�
@H1������W�4��lJ��,���s�����f6g*75j��������Έ*og�3�����~��HEk�a���\��S�^n4��jR�r{��S���Q��z\��cT'Ǩ}��7H���5M�9ц��^�"�ic����� ��i ��f�ϩ�̛�=	��@]C-�=g-�P�GFQ���l�-9����=Ȟ��qD4|4�#JZ)�� � p}G�(�b�4M�T��p�.�N(ug�E����Ҵ��s��5�٭�qE�N6.Vɒ��J�5-�.���\(��K4���;sӦ�'2qN3�oYԶKﹽڙG
�����ch�H%�r'������ݦ�`}��ʒ�0�����J���&�/� >2p����͒*<��zp{��=<9R
�R�~9�Ny��~}��������f{}v��ri�Ui�b*�p.m���*mF�4k10E�U��hf�2�Cm��/"ݖ��@QY���#���3B�w�����m�k�n���f#�"���q�3���W�/�{8u���T�:��t�3<���sڥ�c��]�pތ�f�x�Y�kχ?�g�.g�T̻�Ԍ"�tز���n�R�<Σ9����=u�%F�@��@����pr���*�m���Q���DnΛ��+2�q��s��X4�nN�z�A7X��B�"�m Y�<;��)��-8%+Y�y��w=�O�+��Gm��H��!y�)2�-IA��ȍi3,��xM���MF�X� �eA���Ǫ��������*2�x*�vu+RY����pN��)��*Y��kT3�6�G�+��Rji�U��C
�`��
�RVS�H)��(""��*p���t2�EF�Ӂ�DoWh�w``���$��@�ۼ	�1ߧ��N�/M���d	�'l����>��ϴ�7�A�!�|�A�0�0��@.X�0,��j�3��P�E�kp�P})ߵk�.#O�*�cd� �����H�ϐkw��.R�
���O#���r�H���|�� �x��Bt��MI@�i�*(��n�㔀.��:�9�tkِ�qC��8�u��63n�A�	>�O2 �$��{���X�)����/�����nr���se[M����3!�Ԕ� ��W=%G��ٻn�Ge��� F�d��tI�Ⱥۛ=7e>��#7&��F��f����H'�0��"�q�+�a�5xE,�,9���k���M٪3*s�Vp���.U�ʺF�,�Uω��w��r2���;��K�#��ɼ�uT�`v�8j���(��V#Z��Z�
8��.N��n&�ED}��K�	Ͷ�Թшj�j�����)J�cJ?y�*���	���D�	�F��R`9��1�N+����v�&�۹��\�B1�P���I�IN�F�k�H���q�u{���ɍ����_�[f�F��FF͓�������]Yf1t�F�
&a��z�F��_�r���|��să�5��K7�Bi��|�vc&��[t�ā�[o�U�}�x��\�p���6w!��K���R/�}�ڳ%�"�#�����sx`�Dej����IZ���1V��f8���uf݇dL����ǦC��"q@�1��Dڠ]5|�i
�|JSјp�X}:hE+"HG�� oNC:�-�e ��(���(��MJO!e��Y9/H�l�GǴ��:�b<��
�9Sg��� H@ߵy;�9�h�/YՆ�A.dH)5��QB�����޸	k!@إ�X�Mg.��Gw'��J�7��"�g��^y=��Ԫek-M���}'��@���X� weNNOYpX�5���+/��9�]
��5{p�7��G o��CApT�"5����&�`�hlf��lD�74��o��F�q,�鱎�8Ra+�������^��͐��B�u�`��r`�[�xD�i\?���3�v��u-�H��GD����{�|����E{����P�ii}�r�t^߻�^�O3Y�$o�ݢ�G�#E\��"����{����"��r��q���q��KOnlY�:���iD� ��.]/u��c^��M�������(�cu��.u,����0�	�ފn��ҁ�4�X�W�o��'<3pΨ���.&����c�]���}��V[�� �V�%!�:ƽ��Z�Sz_��~7�r��g�����cq�:8?pZ�6���2�9ʊ�A��!�h�Qj��\����0 ��6�43�z}��C�����l��L^� �U�{��z]�*=�9��.��	���S@BD)eD]q�l�b �ȭ�vb>o�[HP!�|�\��qE��U��4Gm���ښq��9�s�£�~������/�.4eӭ�-č���gձ8���]�-y`� L�<.k�u�|u�ò�"X(��
XW�O�	 �2I=3��.���C�W!%�0�Oh8o�<ض�H���*^Li�܇��9��v�-R�b�e��b�b �X3W��-��'T�9�c�'�����Ϟ�cY�.��m��Qw��-�܆a��X:tW�#�b/�9�s�́\�0�Q4�(��� �68&tk@1���Z#;̽�U�u���	8��6F�M�d_�^�±V'�l���i��Ep)uj-5Z��@�����9�X�7���5ny<�� �/�E-�F�s1�=.,6��*��t a�T�5�1 VMun&HMr6��̵�TN7��a��.�<H����[���֢�N���d�ĶÝ��[hU���5y�����|6�G1�Syd���0�k����ꙑ:+Vӣ���Pt!s�A+{=!��p.�D�ힻ�7��K���MtC�4,u3f�3GE �|��I�qG��{P��D�9�z,�D6��j�9Ϗ��d�]Nn��(
4�L�׍F�4�n�Sݺ"Ru�Ј1�iS�8'��	�ԣ*������X��0�������ij3���V���K��U������H�V��J�3Lx�k�jX�Q�2@&�]��u��t�&OA%�i,u������d�ߠ�<������n!�p�C��Z8,���.lR�Z�]_.[��m�[��0�y܇�0�G5��:��o�~��QD��H�,��Q�<�����"*Ǡ�"x�<�@�ha��嘞R�|.� i&�ڬjqd  �]��ę/<�&����H��2ȵ�lֵ��3T���_2W���Y7m��,���'fm�1���
���������o��f����x�m_���I�R���G�$��5}}e�0hC�;Vvrt����M���z9���1�C�mir=0�<$C!Q��*[���}1�ᢡ���`Pð{�0CGr�{���V�h~������-ׅ�6���R�9��j��<��zZ���u�U�,�w��u����R����P�[[�ܽc#�isb+�qqm2G<?�>-g�#W�"l1�[��"��Gĸ���C9��]z~C,)�s��YH���C�P��p�&bt���L��k��~�x� \�ӈٔ�\ٲm	���2����1֌��=)k��BN�P:�i�
	f�V� ��v�����z��!�2PvC�k�{��B�＠�mD:���I����+x��r/`���/����\�S���Ů��=o���\:��p���5aC_s=�%�LAP���m7 �ɿ�(��zj��6���vGWE�9�5��Y��O iA&���&V��������KD�@l3Ԕĉ�CE#�E	�.�R+�M)�2�2��̆��O�&���C�-$�!�R0��iKy�D��*K���eR�8�J�%_W�J��gp���=e���	h].^Ni�d4B[�nH;����jP*0���`}9�����/sF|���0Gr]rIX��4nu-�;±K�_����(4��.5�*r���pЋ�Eʌ��.�B7@kF�z�أ�x��U����@���t}���zs_�QK�ONy���҄���@�WOd�����5�K)�,���m�k�U����F�������|Q���L^HO�r��C1�bL"����D�b*�5t�	
Y	@Ha��zd�jW�9F�"��V��v��%y������#�����)���
tvU��:wQ�lx��M��B�!p_�z:]x��ԎaN�ˍ��DLB��+Mo3r��µ6ІpQ�wG8�;ɞB;"ȱ����qՀ#�zː=�� 7�V �N�,�y��tZ;��BQ�Q�	��(���q��9��P�;Jui�
��7���δ����)�j3�ݶY�����������8�{<(�����ʏ�8�1�/<"��������7���=k������<����#���;v:���	����b����υ[ܓ�ۋ&�kegZ��f�vߔ�ު�i�|v�W���D6�6�'�2o�g�O�1彇��s�5��:�Sɟw�k�-#�c����qN��a�b����~P��r���҆�Y<��{��M<F���p$�I?�,}/�S��M��x��'2u��DN�e��'\BQ4������	��km�]��yrN}��1u���<^�q�p���r���[���u\��|�:����W�9�~��^7�ϝ�0o�_T?��&��jU����Wz9ׅ�X�5
�p�|"߱ޝ���[�ዚ���ύ�|f᫃yG{�ミ�n��W����ڵ�+���?3��5�ui����7L�ط����-c-��[���Ϗ%zSW�8�aRG�@��Z�&'���_[�|f:��nxa��C
�̛8�9rnd����A8�E���ymd�;w������{������w����A�8�1��w#����m̭$�8�1�q�c���
�1�q�c��8�1��q�c��8�1�q��p��8�1�q�cf���8�1�q�c�0#(�8�1�q�c��A�8�1�q�c��8�
�1�q�c��8�aFP8�q�c��8�13��q�c��8�1�q��c��8�1�q�C��S}���/@    IEND�B`�PK
     ��/Z��d[�  [�  /   images/42ade947-84bd-4266-8f8d-47ba602ec33e.png�PNG

   IHDR  F  p   �pq   	pHYs  �  ����e  
�iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 9.1-c002 79.b7c64ccf9, 2024/07/16-12:39:04        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmlns:stRef="http://ns.adobe.com/xap/1.0/sType/ResourceRef#" xmlns:tiff="http://ns.adobe.com/tiff/1.0/" xmlns:exif="http://ns.adobe.com/exif/1.0/" xmp:CreatorTool="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" xmp:CreateDate="2024-09-25T10:04:27-04:00" xmp:ModifyDate="2024-09-25T10:05:49-04:00" xmp:MetadataDate="2024-09-25T10:05:49-04:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0d4a73ee-b400-4bfb-840e-4582cd31f35a" xmpMM:DocumentID="adobe:docid:photoshop:102aa0f2-64fb-f64e-a33c-390250429f30" xmpMM:OriginalDocumentID="xmp.did:7c2c0979-bd24-4ddc-a181-e94452fe37de" tiff:Orientation="1" tiff:XResolution="1920000/10000" tiff:YResolution="1920000/10000" tiff:ResolutionUnit="2" exif:ColorSpace="65535" exif:PixelXDimension="838" exif:PixelYDimension="624"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7c2c0979-bd24-4ddc-a181-e94452fe37de" stEvt:when="2024-09-25T10:04:27-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d88baee0-672b-48c3-8fc7-826e592b23dd" stEvt:when="2024-09-25T10:05:48-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8569033a-e003-456e-822a-67d8550fecc5" stEvt:when="2024-09-25T10:05:49-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> <rdf:li stEvt:action="converted" stEvt:parameters="from document/vnd.adobe.cpsd+dcx to image/png"/> <rdf:li stEvt:action="derived" stEvt:parameters="converted from document/vnd.adobe.cpsd+dcx to image/png"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0d4a73ee-b400-4bfb-840e-4582cd31f35a" stEvt:when="2024-09-25T10:05:49-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> <xmpMM:DerivedFrom stRef:instanceID="xmp.iid:8569033a-e003-456e-822a-67d8550fecc5" stRef:documentID="xmp.did:7c2c0979-bd24-4ddc-a181-e94452fe37de" stRef:originalDocumentID="xmp.did:7c2c0979-bd24-4ddc-a181-e94452fe37de"/> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��9H  �IDATx���]Wy��N�]�H��%K��U,6���cZ�� !J�R ����.-tb��ɸȒeIV��H#iԧhz��ֳf��hf�}Ι9e�?���)[眵���we.z�BD��k�����R!�B!$�9��W�ut����g�?LS�Zu�VW�B!�BH�S����U���k��&!�B!�D��uA`�(��"B!�BH`A`�J!�B!$�d
!�B!�F�B!������B!�xB!�B#B!�BH�a`D!�B	<�!�B!���!�B!$�00"�B!�F�B!������B!�xB!�B#B!�BH�a`D!�B	<�!�B!���!�B!$�00"�B!�F�B!������B!�xB!�B#B!�BH�a`Y���.�? �ݗ&B�Evƀd����I<���2����!YP7�$ �)=mP&z(I#sH& d��B�4h��6;:�����e�2��G��Ȕ�>�����~�hCi�I���t�Ж)���RӔ%G���3C�������2��G����^)��"��!�<����;]���~kђ)��ZVk�ޓ.d|T��\%��:�����4�O�O(0x��ҥ�#C�*y8ќ%՗��\��g�0G����&G�� ��t�%��M1zh~٠LLU21I�~)�����x4C7A&�2䔒�cJ&5fk�E���db
������~팇�ѫ��z�/��8�2��`�϶��������ӕ�����Oi#�5d�a�^���G�����z,��S21S��ԢA�(�u��M�f_��'�l�q�lM�5C�2f�L锕�]r�ĮQN����X�u(�W/��+�r�$�3I9�k��:eqEwD��[�!.(�P*e��|�lWkq�0b�)9X3�S���"�8"X?\W�����sd�Z����
��B�T\��aUe�Z��1�5!_׺iHh���2���I]�	�����@
_��_G��G��N���6&p"��5U���rP?AF"Na�r�4��.�g��!{��.GH�T({=�C�N��#��\K�������W��B�lW2q��I�hX6�KV�f+�4)
��>��f����l��1.R��eӴ���Q:�;���������B̬U}ÌvY1�Kb	�5���h��ٓ�t� ��Y���J&"U���
ߦ����ܩ<yF�Ù�@���@R�F��N��n�?�� X���f��J&�
Lvq=xu��P�'��: �C�A��&�'e��"�"��Y��:ߖ!�U2��5�C�ɐ�屶�J��oq�V�=E{��q�O���͆������~�L���Ի]�"�����P�A�ni�ܽ�U~S] �+rޛ�閔x�,!.���pF�`@�湭r�Z�x72����������B��HA��v��,K�nR���+��xӜV)͉�n�9\���Zى��\���)��������y˂-�O�.��֛�\�,N��VA.T�W2��i�k.��N���F���m�za�f�
��Ļ�T�=�ZdCU��H�'�mW5���g�
�3����r�2@���������K:#��CEr�>�YZ8pF��'�딣�F�j���� �:�o�����!�ik�u�F���E��#�h��õE9��(���v"�$�g���)��z%??\����!{�(	�A�V^��A��Bޢ�"'	6�I�@~z�(�ˤ|`�Ym��%�z*G2���U�d��.���b��-h�uq��v$(�Oo�׎��K�@[�;�3��<�n$ΰ��Jv�^��g+ݤ�"=ɺi��M�tӪ�A��L9�<�Cوd$�F��lݔ��k��DM�r���ZLȋ]{�X���I�݀~
�<��!HL6H�~fc��X<|�H��cA&Z`��a����*)a�%z�׏�إedIzv��g�?g����*��2��)�=m����}a|�ko�0Yk1�ll����+����"kp'֢�Gz;���M�7��;�J�~kO��lNYQI�w-m���)y�W�#i�C��@��컕<��uhQ�������Q~u�P~|0FS�\~I9�c���M�mz=���<��!2A {}P�i�ms����*�:J�tS��D�Z�V���!C-'�tAy�|S�Eg@&v��OK��a��!������.-��OQ[�O���+{�T@�O�����+[�d2��b�ebl�m�����҅�o�^�4��wlv���b�����������iL�@5%�.��<R�`dWIfa�dT�*0~}���zAzZ�I_GcD�ZX>��A~���T/�#����t.R�T�����ȯ�
6P�}���k�|V;$��і���Nz�TO�IU�\�d�!�p�dMV�0Q2�˵��@o[����W�p:����Z�&��*MiG{ꠛ0�9R�uS��M��n*�;W꦳j].E�oa���\Ӡ+G�;�ں	�OT�!#�L� J6����8�Z&�n:��&�D�V�#�*��#S�e������IV�c�'�u)�+��L�]T��^�H��eM�Ȃ��O�T젟�i���U�2��>���H@r�s��L�r� 9�df4��f_���z-$����N-�Q6�L��O%R.0Z2�K�j�������.�-Y�ӣ����P]�S��Xwc�t�W��m8`����)uc��{��<ۑ]6K��gic-P��%Ӕ��&ySE+������P��UF�V7ʷ����A���V'P�Ȯ���b��4EG\9�+�QkpB��q����[_/���L���j`��_�iu��	��ʕn*��nj�M�"�Mh�@��OR���i�a[/����9Z?E䀏 I�l\j-AϥSZ7!�d�?��A��2y-�D"���8�9�	����֑���̂	��I�uǇ���c9�h}ř0_�Q&�&�=������h��^�R�����X�p hC����):Y�/�L���f�'T��:נ��e���LDb�1��`�/�оȔ
�0�	��H�A s&-RQuE��}<\yy+$w�R�xH:��eK/��#\�b�(l^E�-r*�굀S+t�D]��X���Uw4��G�ތ�����<D���g��� [�E�HK�Rk;O_=M��u����{��@}\����r�>06UX>���"�MX����2��ʔnZ6��^�BqǼA݄�v*���������bə�0z'�$�p������]Y�D�O���2�J��`(dbJ�S39)٘�Ndn�U�B2����Տ�m�۞Z�Q4-[Z�k{;;�+�ʝ�DىC�U�^�=?3]�ɚ�
��M��#��s�~��������ԥd"��FR�o����O�24&e#�X?��1lP��]ޔ�1U�#�Õ[�DG�g��͂ܦ�4N"�i�dg1q,���Kޔ�c� ��#o�j]�8�G���@��K�Π�;�NDi�@9��$k(;�UwD��n哛h�þ�ϿT.�)p &���~�E9Œ[u�d'B7�V�7�nB�t&���.j�((�����-h�V/6�A��^{`���?o�����o��9,Y>(��k�r�����F��*���J����E\�uy�^ty�Vk��L���^wWo�>o'��z�"	�� ��Gƅ���6�*�LQ�����ޓ�QE^�����/�	8��mc �j��u��������^�L�}��B�kE��p:��'
(��97h������7Icg�>[į 0��/2rK�B?r�@�-b�;t��	�����/n��Nh�nB��8~y�V�H�tS��n��M�@���J7ue�>3�V(T���#�7m�n%M:iP\%�w�ʅ	���ŪF�܋�����,&�N�z�:���p��������4�?C�I����w5]6�_n���{��lw������W�FcW����j���t͔p6�X���&�f�����_����V�l���"�xO���)K0�h�k?��s@��L߶K`���Wxg�Я�?c�v�2-�X������}�	��낌8Z���8�hJ4�
�y�t��%]�����n�\x��'�)���5��Y��u����K�-�s�n��p��%_dHVt� ��XC����@�{��@�b^�
I�d(���ר�������Mfb�J�$&�*�N$�^�`l�w��9���˛���߄��[�Z@e�f'�mGr�p���f��[�M 1[�}%�g|�l�%�����8�̱�p��V�gy�?��D_N���e�Zٚ@��`�&�$d?��0M���s�9B߬��W֭�Px�+��	K6yU+�hW�
F��,}��x���̺V�d2��nR����.�ç���[M��]<�����Y���t���]����[�?�-�~����pI��cK2�s �l�ݮ��@���l9v�퍐g�1�p��$�^W��k���'�~��5��'�1h�̷�f������n��`�Z����k������Y�p����s?Q4�Z�������u������'Ц���\F[a�z�p�l Y��9�I[��g�`�X�i�z��h�n��T�����-2��.��%��j��a�d)�}]�2�#�M���M8��	g��	���F�;Q8�u	k�3�]�Ah	D��O�H��s�w�
��"[ȟ�V������?�%~�d��5{�eLb^���Π/ێ=g�����n	�3�f�9褅R�g<l�
��)����
����.�>�-�:k��a��u���3���n$n�Ѯg���E�1b���p���hMP���&��,��8tp�Z?�����s�L��)(r������p��T�{5������d���atS�S�@7)9m�~Ƹ�⦙��i�O�����0�\��	��m	�t���k����Ɵ�3������^�z�Fգmʦ��N�@o���nAy�>�����p�'h{�ጣ�s�Fk�"���^?c��	?��/Mqd����ZX9`B$v7*����U���U���P|�6����(Y��c#N�nˑ'���n�ɂ�Fw�o�,���P����xy3�r�%��+�n���rG+�[xL��8c��
�a*���@���}���v��0<�
W6Kl$-3G�kˑ��t���[|����M�~��Қ0���z������K����v���M�'c��=kU�ڔ��s�֡&T��^Ъ��@@��og�K'Nnu���C����ۮ$�hc|�BsǓ-���|<��p.��N��}>�3���N��t!}���J荾SWK{�+���y.���n��h�8��z�9�i,d��Ї��6^�������V�<����Nc��h#3��^�OEwm�������aw������`"&�u��p�>���	�G�B/��H��O[=�[	�Xo[�q_*���'�߮��H�쵞�haV<�A�]W+\��C?���3���D����k�����s܃��TM�k��^�7��N(�yK�p�h�6���h�����(Q`?�A0��i6Ѣ�j9g̒�*f{`t�Ǚ �9��!_)~ �FQ�Z�nUk�v:Q����:��<[+v��Z�;e�1���	]��bE�~a��n�<`/Z��MBl��t����9?�7u������0$��Y���� �O꒫<��@����vp�:QL<��_WZ��VO{]����G�k��_�O��^txx��
y��X��B~�7�>���~;�ė���T=�1��2�2����<�,�q�lh�4��1X��;�
2�m5�Ӡ6Vu��ʹ6�D�fy��˭��B
��(��4�;�x�6F޺i�u}�^�&�u@��j��vX��p�4�sr���Q
��r�_?�����K&�N�ɝ���K'�C�^�yf������+��Z�vƼ���	��k�ވ���CEr�ҽ�7��م�w��U:C��L�ll6�8�V<ӄ!�qV·������<쭰50��#(�YhQ��"cloo�{�
��O�g�^7�#8��X�Fn�bc`�ȿ��0p��<5�%O��� 	&��v�q�>�����z�v��:a�'r&]�O�w;{�Lר ���WyL+������S�]�{mk`t�4�L`2��T�כY?�8E:�g��\����J?�#�&�����&|m�2?P� �4�7?�$g�90�QA����m��ď�u��S���|�M�)���b �l��B<v�Plc���MH�#<l ��u���I�Q�xO~{�;��s�>d���hC�9(�c��g��A7Ђ�y�k&��'y�N��L����ٳ10��aJ�!a��P�/�lİ^={�<b��6����lV�8�ҏ� 5�u7�p����]�d�]{����l���Y7&=B0B��:F������n9�`O?���`���C�z���m�Qn�n{5�_�T�+�hr�tO��K7y���i����G�'������=�aX�%���	���W��kx϶Fʺu��T����j�����6-�R�'�}��{�e¿6���620���e:n�*�U�J�G`�|b�u����2�vO�	G�z�.��3hS`�b���W����^k�^~���[�EgU�0��m�~E�&C`����F�=�E�O��'Λ��i�������@$�LGj�9�-�Ȅ)0�z�����)����������-W2a[`��K?Yz�L$`�**^n�TL��l���:���U`���� ,?G��@�hG��	���,��e��|-Գd2zz-ܧz'8�J�Ff�_;� �x�t]<��=�,���Һ��J?K8�r$K*�s��ezV�6�~�xSVv�z�6F�=��v8�g��g	�G��wN:�b�{�e��}����;�������c�;�'?'����f_��{���=��'����dU�V�r2���,:Gg�a-�F�l��A����:GW��3��87�ɘ����'�y�vF^�	A����䦛�B� �ƒ3CPM4��Y�2�a��ڕ@C���̢Ԑ	���S��������u�������N����o>.(����Vrm
� �10�=��������ˣs�M�t�kK`��b:L4���#���F`fq�k1�����X�̂I28�}�U�UbŜh`xM�	'����Jͺ��s�<t�-���L�_&pn���M2LmtB�
k�cgy<���iڂ��"�:C��сt�꧄�i�z����N�d"���U���!w#Ӈ�m܀�3��o^�%3�LR�������!0�jZ���H�uP�<#���	��y�i?�cm�M^�EF�؉<w��L�)�r֒��Lk��J6��V�F?��Z@?uK�����m	���I=G���F;O6��pءA#�tvH��w떃����<��	�Z����<;���L���1�7'0?�_�����;�������Y���M���<�)�#�qG��� #�ȵR��H��-���[���{����?�"�4BJ���]�i�zSg���Js�� ����(͵c-L�#=ۮ)a���@��y=�"8G�4�4׬�IO��><G��g�$ǎ��W�" ��-0*˱_&@z �Uk���e��Œ�,�����[����d[�{P�Z<#�OUq�S����@��4�!���k�0x^�Cz
��K�K`d�:�B�Z����0`�Z�{�D�z�!��M��o���:�v"O=��!-06;��S$�&0���P�)�����^���y������d��Ggx���D���1��<��=�a@��l�S7%�3�R2�a~/��D��5�\tJ�#�Z�e�q*����0��ʲD&�#���p��j�86鯴ѥ�I�⫉%-�K���
cE���X<���G��l�21����Mcg�%�/V��74�bmy����x�|�z�3`Ǟ�X0��^�����3����@3�_0����`-<�?����^z��x�<��TZ�<ر��)d#��)[֢'(2�b��H�u ����;�$��7�Q�G��@�]ۍ��>���;z�iQ����/;��-��'�����h�x���'���:z�0x^k�����齴�ر`P6G�T�^��n�Lt�z�D@��%6�{-���X~g��~����^������v�D8|5{L���i�T�m"�i�GS���H���뙲a-�T��ڝ.�.�0ϐ�}@��d����M���M�d#<���.�DO*�k����Ж���Z=Ky���`'�g�|�L��O!����Ŕ�󆮾�I��Z]7���h<ע�9%���4?S����E�:��T��ox/}�m7vڱ^��ߕ*�	�����nRz���Uҳ��xɷ-k�m�[%U�7������.��R�;^2Qo�Z�F]�c�Mk��Ц���7��9�C��:%�zg��Y*ﵸ$R6S���Z�ڱx�KzF}e��8�B?O.��<���n���n�M�tJF� �,Y8Ag�ZT��v�*�ά������~<K�3����^ح9�.6[=G��sR@?u�o���W�� ��OqS�m��
����w�ٞ�:ٜe�^_��=���v�3u�Ŏ����h�^o�E��y`cgr<���D�=6��2��`�ޖ����M}��ɞ��ғЯY%���t,��>;�S <n�785#�D�Lo��D*���j��w���6�m��#E��R',��p���D��KY���@�������J�3x&�]���ޡlg�^(Z��0�����������h�O����L�����Y�g�Lm�K�U�YY0��9�Rf�$�3=-^�ɞ�8�d~-^ϓ_�{0M߲O&�d}��	l9�����^W[$m=�R���iEn����0���}�����Ǟ}-^�������g�tlu#��p�>[���h{�N�:0B{�hnQ�-���F�����9�W��M���C�z��i�=�g��x�޻M๸֐	���s`��]W����6U)0!�<�v�W�Y?���Mv%�y�J觜��Ϙt,�8h�~:���-0������8Xo�L��p;<%l��Z4�'��U`�����w_:%ySW�_�t���=�{��o������Ɠ����7��=�Aў9��rt�Y��Kj|�?������b{�uey/���T�R�Jw�Y7�h���*�p�@��	?F�i{-���5tfHy��
��zPOn�����n�`�L(9�e���0m'|yɄm��!��Փ;GO=Ox��}�G�'S�Cj���^�*0������z;���o�����b����*V^���J��2�q:2�=-g]��ݗ�޷]k�C���hy�i`�]o����k��eA�h݄Q�ݍ5�lm��M;���B_���ia]��N�Z���Կ��@C�}�v��p��I^�
�#x�&���rue7'��^���m%~^�ؗ��µ��t����>��d�s����
���3����?������a��;��l[#����M3܍^W�aɟ�N�FW����~�l9�b�mgs����[0a0���I��z�:@�^�[`�\�10��`�_�d�}��ؐΜ�:��S���	�ox馭g��F�*�i
���Jn�U��߂ği*�t�m�گ�{��k�o��ז�k��JVa��]:��-�헇�
y6a�Lx�������%ͮ�*���W5�W��A㷟�����j́QwC��T̗��r��>ye=^�p-���Syr�t��-]�.0�p`pޯpƏ4��H����w(���F�&�U����c���|��M��t]8�u��ٳ7*�k��Ľ�i�ٳ�+0�*���$�j���N�x�T��T�d���ʙ0�W]���\�~�R�@��sJw���W���A��~'�������]`�ѸO�(�7�r���y~�`)2͞I$^t��g<������v�p,�p�(w��'�����0qX������g�3b
��觾e���x����Ъ�T����4�sJ7���C�yV�^��Lz�|�N�@o޳�Er]Z}�{��Z��OK�r8�KM������zZ���ܫ�H
B7����S���^c@�i+��+�}��Ȱ	�6o��90���$Ԯ���߷�f��]`�8�o�p�eǙW}1��t�m�w������z�������.��L�'��]_�9��5��	�

��WU�;��gwKV�_��t��j���J�`
���[��{���*�UɆnB��V������{��w3��$�`���Yw���O��-p��*��ǌC&
�� ��v��3f��}6��v�����fW����	�&�>m�	��5�M6{���U���2q�=��d�	_F8i��s�}���Y��|�_:jw���������]	7*)W���3;��Qau��T�O��Y6[��8�����"�^�C
fn�A�Ի~Um��8d�)���a��$���F���CZ����_�Ǐ*�.�Y�-�wH��7X]���-�}p ���D�_)[��e����u�Gn���v���*���>�	��@�h��^�f�^��[�à��ӻ��G��>�ӂ����W��6�n�2z��������nدQ<z�P�����*:Nm���"k�����Hb??\hu{D(�s�H��`8yz`@�O�,��n��t7�����c�/�/�ޞ=e.�cLqgn���l#h��<�������$�y�ykn������t>�O�l<S@����Mh��kŞT7�`���&�3֋��E��� ����_7��\�t�i�:���bkh���}hg�u��H~���OU4���c��r�Í����9R$~ ��)7�0��S�fۛ0�>�������=s��"`��M]�������|��W�N�$�so��,��^���k{)8T����7N�ȉ-V�7j�٢���@Ⱦ:�F����"�fr�1C��Lzf�u��n?���g~z��\R��'������C7�+�T�u�]�t����M��>Q���[�G�N�4�! O�̵nl4Z�a�����b]��?U��S�����Z�'ۆŠm�k�W�Z�G|���+{�@��&{�8d���o��eBP��_� ��P��O�F��O�ɩ�k;�D�W/�d�G�����zb�����Eڎ?/�6Iz��{(�6����C��M���ӵ�Ϫ ���Ц���I��������ux�rs%�y��r /�h�\x�ˣ�r�gSm��X�t��I�c����u��M�$n����^/~�S�������8-]�,Ơ�"�l�~��q.W;�~믫��~b`H&��&8����?��� @&�*�Ti����Fm5/*{}��^��>��m��󝚕����b�_+�6�_���-	M���h��uXU$�:0��W,sK��$�=�F���سR0cC�GG�)����{JH�]��	�=�i��{����՗����Z����,H���,�vxM�����ѫ&0�{~Y�q�:h?�]z�%g�"I&�L���:���)�f�����y��IQ�I75�Ì���J7����*][��?݄��p>L-u�Cp�^ț�F�I_{��M[��H�������<��*x��:�:�muЁM�^ 8}��#5L�����u�Z�?h��T{��%m'_�I4/�[�Dw���5�u�lS�w�W�)w�bI&h��~���U�����F���ݥ�7ט���UZ�>%���&�#��S�xnR���S�H�r�}值���g�rD���5I9�������Ƃ(�=��B7�o�)������!��e���"�7&h��Op ����}8�P7��>��K7�(���Z��I�
݈��k�@덟Z�F����E��~~�U_�b�Vm'��a�3Y��3��L5tڷ�#R���D���z)6$��Q���Z����g�$��9  ���W�7TX���^�����Q���۵����>�����9�~Z�a���^`-�10���H�-.���_������z!G+�?[f�0���l��'j"��gv�L�xph�F�V��ɛ��"2��;yY�^[$�8@pꇩ[^<��T�nC�L�7�Q�a��P�V-���)	y]z���W�f���v���v�:�`���ξ�^H���M9�a���Mպ}.�nڥ�÷��_7}S����>Ynhox.[�^ۈD��"#�DE8G`v_�0E�k;K=���x�V��"#71�Z��x��fϟ�{���;�96h�o��a��`�7� 5w�҄��H��o�{��w �V6����f��SV�#8��a$w��]er��6�D`P���엷.����BK�<g₸�d::/���������ycY�����,�2��s�Z�s�����פ-���vF��j��R&_�`l3�Lڎ=�+�(ӧ�ħ��E��ty�ʿ�����P����E�t�1��	��	q�MJ��U��k)���^ ^�ԁ��nڭ��"�`b�^�7a- �@�Kt�X��n��9]�8�;��rԕ��VN���:@����A���](���t_�DS�P�k�DV�Q�d"{�I�~�������Q.{M��嚃��N�O}Nw`-�g�{����%�~|�E�F g%�	�0���8�h��G��U��9$�k�`(��e�d������j1��f��L� `�J,[�j�D!dX"�3��U;��Y�^.��^Ө��^ a���S1G2�+b�P��Rw��	[� (��w��cGu�[�G�zpZ馋G�t���&��`-z�SG7aoſB&�6�^s�Sު.�����o,��A't-DZ{�^�	Κ�$8:��tH�������͘�^e �T� *ذקZR�u�퍰�7�g����܌��wR2[{}|��5B{����ڛ:��l�T��L>�l���06[��O�1��G�v8@���M��Z�-����p���m�QB�6z��a�K�#t��E	��M�#y�L�|u����&���Q�w���`dv{�˺�!�d��ZL�*C!F�����\��(�)*~�0�6����r���K2�p�H(�Z��0��⩺\�Y`P�=ʡDe6��������L\HE��A7=�,�ԪeA�Øu������Γ��JM݄�>��B�D������$q�g�)Q�������&u��S��S�3������V]2)q�~G�WfQ�~*�u��fP?�z�~��KY���B{jT�F�V~��;�Eb�땽��OJ&����DsV�@����):{�D�OR�^$4�~Z�(s#�كIM�i���LD;�g�6���#M"%�#��?2;�]�$�"�R���9��=�8 6M9"�ئ���}JP��=�����j���F���L���G��`��9��9}���� ���!��L�����Ȓ��t����;�8��da��X@�hs�: cL?��B���S;"�8�p��(݌�b=Z��L<p��{�u_>� N`�`#36�����,��!y(��n�L�C��A���Pݤ䡷cl�	���,�u���N�÷ȝ�"KfA�t]<�/���T�GzN�Ԑ������7Ek�Pz�	N���{qcpxG��*He�T}��A����
`��i�,�~�l�'G&�)Ta�{��:��@(��砟�$�A�Ib8�Og�e���I�{-�^���^�r��k�'(��$��Eh�ճ��J��(�l��/�f��Xl6��@���R��{GC@�~��	�Ͳ�*�E�â#�8�.L���Tk��vP��ZDj��<Ǫ@Á��1���GGKo��,�Q�^S݀�C)�LR4���R�-jݴ�)��E(��Mp�!;�G7a<d�]J&�#L�i���� �V'� ��*;���q�
���R!o[�,�ύ��	��=�.}OɄ�'2F�����T�zA�=���r�!5�� A��}�T7�����9�6�Y���N���Tp��a�ϟ.j�8C/�	���}w6N,@y�e�?]ؒ�i�W�j�vAS����A �+�s�cZS~��a���y���P��}�C�CY�u?�]}��MHR�*�V唿>̞�x������l�X�� �I�o<�s��8Ӛ�n�+H~��
]M��E�W;c	��G�:�� ݼo�f���\�]�mvQʵ΍$������{]�<�M2�[G����Bt��l(�"�F�x�<l��lyq�%S���L��ҩ��%�u@P��~��N�v;D$�@^���A7�JF��M�T��h�u��ȇ���L���D���.�ɚ���������B��2�M�늼�&��A?mPW�	��-g�~�1	�z󐽾`{�c��Ƀ6;�It:���� ����og��2�];����nU
�߁�`;#�c���8{ k���`���X��m	�#l|ƅv��g����5^P5�DW�����6��Js����2r�'�9��/m/��J^�d"�V�hA�2񤺂�6)O��k�^�Ɍ��&d�T��^>ˀ(%���m�^w�5�{��N��^��`׺)�6{Ʉ����f?@����u�8\�/d�񀡥(+#6��l���@ @� �=h��8�C���c���^9d��ؾ)�X��UңA����	�ԕ.;���$�kLx�	???\��uZ7uȪ�]1K�M��M� ����}�A�&dj��(K�@��mC�	��Ը�L����j-��f����m?7����!f��jl�X5h����^�q���@��Ft���=���م��٘�6�mg�����d�ӕB�b0 �2S�9�I0pP��=Ґ�?C�%��9���~YR�-�Z�\<��W
��A�AF5����@�k$r��U|�+�d^Y���F�tѢ��1K(�8���1�>覥C�i��M=J7���Z��j�����P�8m��0�U��j-�~:M�H$A��t9ْ��f��L�Ul ŧ��Ttp���eݲH�ż!����^�#G1������ z�dDEl3��0;J{����C&��h���e\8jdڐ͞�l6�����٨U6����������!?k@k(��ק�gN��N|�`�T9��&��g딋�h{�98��"�
k�u�fv;`�p=Q3�w˘�Ò�>e�t�J-��=i�����L_,�s�L�+tS�T��ky�nJx����ӗlD�Z8�9�	����c�R�� 6��ig�:��yu��g��H%�	�'�"�Q2Ѧ�ӥ��S ��؂`���O�k�E���F�N#�5�Fc�|\O��Z�ĺ��%Mj�,�fun���k���cP�T���72K��p'$ڙ]��B��;�ŝ�lh�� I ��AϟB!�xB!�B#B!�BH�a`D!�B	<�!�B!���!�B!$�00"�B!�F�B!������B!�xB!�B#�4�~�>yvw�<��<�뤐��_�Q��k��$~��D��+g�]�ʼ�er��U��B?�{��Y8Y���o$h00"I�� G�TFׁ������n�x^�j����w�ǿ���9v1n���-�o�v��+���?�Y6�u�#��X��3Q>~�ZY5oRT������J�;y9��OCK�<��I�!r9ѰVD�ς
#b�g����M�嵓���G�p$�Y���ݿ�U���~��_������]+��%UtB��8�u�C^s�9"=u���� {�w�5�B>����L.+�����?��գ�=����k��g��R\�A U�%�&��	��֣��O�5���Ӎ���Ӵ� �p熹�Q�/
��к�(�"�NS[�(C����.2��%|���jm�bՖ��w,�Ȑ���T�vӢ+�VV�U��ܾn�(=���ۿ�G�0J�ĹEp���3�Χ�[�e��r�����=��h��
We���*��o;�.�$�p׵����DA0IrY��{
'[���l*��t�<���q9o0������y�:��F����o2�za���]e��r�(x�mK�����y&�>��W�T.v9���tV��⾸?��3��>w$�8����`� ��z��7,�橻 W���I� ���������~n�[���m���(���ֱ8oP��gͨ�<��d4���{�FE;�^�W�3�<B�E���ᙆV�7F *?��N�;��p8�^��"���U���5U��9# �@��������u���t��w&	⋳�.TF۰��^~�JM�}+F�'��yٶ�Z�~�� Y�ķ�י�� >o��j�=�P�`G�����<�K�;����-�-���?z栧���[�\�v��o?�m�����30� |n��4*E��������~S�0!�q��v�"ړ0�E�zoQ:�/U{~~����k��5�d��Jc��W&�G��h��b'P��B#d�F��G��=��6�փ����Q��i��_�޳�!�VFf��|�1P ��op.B�n��R6�=ҁGPڞ�v�T�Β�5NϢ���H��ΝR2�g��g��.��Y0�L�7H�8�8��H�D��Y��U�ݱR�:��t�� �_�x����	��*�A'���7~��Q�N�2�Ⱥ�<v`��EE;>O� :-�/�:���������A�j��|�h5����t'8!�pqơ�P�p���9-0�E���S��v�4� Pu����/P�u�?��1�Z�J�T�pq�W�xmCp�>��a`D|Ch��4���u\�ja![���I{�31r�J�;�=d�#�"����O>88�m��@�6t���5����82�A�	�\�x9h!
#�M��w*xA>�%0,�:f�	H�>�9��}d���ݸ�"#q��p��J_2rh�u˦�j!BV�i�c���p�ё�͜3w�zzG)e���w���r	�}�Lc؟�y��+�~�d��@ː���H��F��Q�Oh.�
j$��ᜣ��&l:ۼ�`b��U.t��9���u���sd젵a�hV��!���)Hl��B��HZݠ{BA��3��e������RJ�Ohki$�h���f�-��q;ǋ�P�``DR�ںV휄;x�D2���򱷬q�~�i]d|�󷟹U��qd��$$B�GO{W�Ж����fB[Kc}��N;]�~2�O�F��8c)�zm����	�^�I�y�X�~���5
��V�m;B'����7rѫaԍW]���VF&��#��XW&�D�}a���9���8m.660B�~���{����RB�nWJ��-�v�83jd�����:������?y�3v*�9^�`4�� �{�z����kX�ϯ���J�6��I���)7&���er3<���[F�
=��y�G`�Ѝ��?Dr�3K˱c�|�΁�#�J;����.� '����N����<���"��v��������)�L�r�>5� 64Yv L�
�PĺE,� A�pۧ~!$v���O��p�΋���q�Q�60"�⇟|Ө�ܡ�V�(�����1� �_�p䊽,nc��N��b�DVL� ?;8]��p�'�p�FX��v�H��	:؃r�����FU6�}�r
�dn��qǡI6Q��1��P��[`:�v��r|wd00"V��.cu(� �8 ����K����8��J��+z���ZQ�}]�Ap��ZS���X�������<�]����}a_��������!��|L��8/[ްf�9*~n��o�{�װ_{�U!f�=@�����֍DG�9��_��H�/܏d&��Q,ϵ���������sG��G��P|����wlpmS�t4~{'>t�J�vE	?�@��[��Oݷn����1�%�}�Z�N(��� ����z�����y^n��s�����ў�!tP��������κ�����E��b��G����������Bl`+ �x�x���Au�FB7X�p��{۲�<�p�qxe����.o���˷�O��]���9������̞?e��w�+����X��?��|���¶ja|�InB��a����F ƞ�묡����2	�i�6�Y�9�~$�����Sv�'Dޱ::�A�	6�zM�au(1������3�Gw��a���������فCO���o/p�M/>c��r8ܦ�3t�4�a�c�66����u�G�$��|�3���D��a�@`@9��=}E+���4Z�
m�� ��n`�~�)��Fc`�(�= d4��HXJ�c�v�Ɔ"���T���}�98���Z�sp&����F`�wډ�5�����&:x�:��*ݘ�czt *�����_�e#��� �6�d`D�`�(��s��ZV��G��X�y��Q>~�Z�2?{A����E����#Љ�?�#��mEby|����)*�;7�ʧi@ ��$1D2�!�00�V��>C�6�#�xI�mt,���Ѻp*�h����)d0�9���unS��q�ƹ����F_*9��$���ޱ�U�8�=l)���}�	Y:����'��$Y~��!y��W��>�g��o�S�{r?[�-`��� ���l\�VV��Ã_~B��YN.��	!~�u˦y�J���:Y:�BW��o�q��u�2#�N�gV�B�gCUy�L*͓��^9rfp�3�����ۖ����Gї"6��h�*Q<6EB!d|`0*�'�x�����ΞV액=;��8n��"��`��3�5^=�R�O*�Ӹ�
s��[��g8��Ue,��%�$�YF^���{�|�&)	���``$�%��L�+������q�����4�'���bB�za�xtP��b'�����a\S���p������|���������Q��������֔{oXU&����C��۽�HBb����[7*�	�}�\���kљ�P�Tyq�\5��߅�� ��=Kǐ���������a	FH��]T�$��d�=�#ق
�p�ӏM�M/�!�ؠ5�-�Q%2�H���������?���'h�cO`#Ӄt�*}��H�穝'b~O/eA�qS�p<�8';���߉}z���y0NIo��f6B(v�uI>���[�&c �LD��_�a��c�4&�)�h��C`#b�n�������U�Ѷ��,�<8�e�pf~��S��F e�N�.�բMK��}�AQ(8K/48B;ҿ302�=w�@{?B4o���)��:����y��:��?�V��p?~�Z���B��;7�vܚںb�"8������=LA=ؒ������(m��8�}�=�{��"d�0*�޵Q�}ռI:뻇U#BH�,�Q>��Ƿ��q?�L�e`Dl��:�60��d�\��eS����腘9��]���J 뻇�!$J�*.��ᬱ�s��
���2�:�!��3���%��!�2�������޸��hW�AB	��AmC�v�p?���x�FJub�P�����V���s~$1C{_B��d�b�F��9玔E�!�8ī���w��H$��Ώľ��<{��/"��:�00"�;Ț��=���BH0������:�00������Ã�����X�M���ʂ�p]� ^�ZYa0����J��D���Q��	�zwp"�3Ye��b�%kV�9^Y�T�m$Ɂ�`'\{p�:*�#��bL�����*Q�����H�hh�v:6,��i �"$���%�d�� ����:��!��,�	��N׵��}7.�i`�ސ�9?��������$��'�����_3yB���F!ޜ�oΘ�zDgh[ick0m8(v�u���7�k�T�?/�Q.���������h�]�W�2v�l��]+��*V�b�u|a`D�Ύ�{�|]���wl��?�ظ�������a�a�u�v6 �k+ezB��jD7(v�u���
mmt�Op�T5��@��S�����޶l�iw@���>�*Q����/�HҀ ���v�������-_z�1mrF�������t���b�a:U�s� ��n�?�츕-Ϊ=���;�;��>�/��uÁ���K��g����FU�s���M�ǫJ�Cacy����7�HR��2fKgOv �_��M�Y@KC$�;d�޸f�nu	5r��}�'ۅD��_��;7���z@َ5�C��{�^q�9@o(v�u���=�_�w���_�z`�*�g���/�&�}��7��ڸ�6/V��ǫJ��c�c~���:~00"Id: ԡYT(.@(Xd���+��Z��8Oʋr�υf7B�����v��9
>��e����=�J�[�Ӱ�3)�o��� �ʂ�p]��KsG�|莕W�8��g��皆�@P����9�%������$��@�}��ruFܾ?����������K���,��ϸn_7;"E;���
%K0r(v�u�dŷ:?*�}�tdC,0���s�E�G�^%�ް�U�$C{a�>�!65�,�5s"r.F��ؖj�q�u��S�p={m*�P}�i�QĚ���	[�"��`'\��z�m��0�ޫ:s�;q^��!:P%rK���^<V��u|l`�v�I>����EJ�=�;�'YW�� �C�4����=�.��btq$쯩�N�3�N�d�nP�,�	��.�F����w���,���z��X&�dE�ul	l`D���=l3I*�� ���e��~YXfbce�N�.$h�E ���$�������	@B!�~h��O`��|'��?�w!�B!�60"�[������m!\B.�2!6���B���nZ�O2�&�G_<�q���u�LLc9$��00"ց�*���)J�d�B��3���Pņ�N9u�Ev9Oǅ�<�Ρ�}�jyvw-'�Y ��pxe�``D��=�/�E��eRi������ ��������X�Vp(��C�L8�3��r�ƹ�qy|�q��D�o?w��-��@���y�u�d��:z�ϴp]!���z~�q��s��A�a��aϼz�AR�H�AfM����_nZ9�'pGA���$��虃�R�n���k��ҕx�.��y�Q48�pZ���ĉv���$E��oݨ�FS[�4�v��Ӎa�1oj٨��w��Y!��T�6�u�'�jeKW���ɗ~��B��}莕�
Q� Ƀ|?����L�H��Adp$B�)�P<��zLN��7��%�.���}q�GEE��f!��9�8mKgU�����+�p]�m?��|��U�ۯ�u�õ�r�L��� ��*/U��Ą2��A�2<wn�;�X`��x3�]\�U(ܟ#w��{�� ��:-��H~�J�0?�.$�p/�= A��[�\�����<�+l;\h���_޵���X.�H̡P�g� �_�p$f���dO1
�w�;_|��Y8Y��QqE��q�ö��9����O\��p/�=`O��g�X��c��TI�z��O��-g
�}�F���m� ���$G�B�c]с�x�m�tňʜ������������6 �-������ÿG�ׅ�P-
��'����z�0/[���N�����$�G0�!���d�����p ���@�t!;H�ׅ�xl`32�S��J� A��*G�"1q���$��NSI�}	���}/�cw����t��+�q���$�IU�]�k��̂ie�~╚���s:�58�00"I�"8��Y��x[��q>�U�"�F�!$`<�[���u!�Ă��ˉ�XWtp?'0*/ʕ ���$��3M��˧�_'�:b�!=��_�CHP���B�ׅ�-�~����.����H�xx���H����O�&B���͋�.v��CH��~��M3:ݐ��N�I,\B��H�@�܏�98<�Fl#�A�gM�4wtK͹f�6;��̚\,�y�2gJɨ�}�1�<���*طr׵�F������:%�|��#�ׅB�	#�T�1�Np�}G�ݐ�����TÙtv��iƩ�N���
M\BH"�A�%^�n�7A��I:^�jЛ�c!�������� )�W?t��{�B$�!$@�8�R�Gj#��T��:����gb�3�v�Բ��$CGO7ʣ[��:GR왻i�ϟa"�p]ϗ~��{�0��aw��a�莍sc!A�p��U�#b�#m��څ�Ɵ7�?"���6$z���K��'{P�*Db�$���!��9b�.���F�����K��m>(w*]�?����/�f����!������	=E�ďx�G��3��;ʙU���u!d�Ɩ���h~U�Ē�����N+#/������>l3�����c������4��H�U�10"��$�����8��
��.�\�pm�p� CFb���f�m�ě�<�K�V�����7���j��R�=JoX3늭H�`�vPa`D!I���f"�p]�̓;O�p����>x����6����Oh{�s{O�����-��oݰ��_�j������c���Ͻ7,��cN���B�E����ݵ���U{ຐ��*�Σ����op�Ϳ~�Gs��+Z�9�m�/>xݨaUh{���M�뉤�����a~��!�X �g^=�M��u!�2h���}��R 8������mǣj)E&��������{��G�N�m��p�d������s�#BI:����BXׅ�+������]��g���B�c�;�z���W��iԃ&����Q���T���5p$.�KfM�G�G�{f�G�JBH��Q��!�q����e���)h���vT����.Vec@�mp�q�a`D!�B"�����ۖʦ��<�7z��Ә�F��#B!�f��h�Z�p�̝R�y 2�C��5ɮ���E���!�B3#[��~�d_�5��?���B!��Q ~��!�B!$�00"�B!�F�B!������B!�xB!�B#B!�BH�a`D!�B	<�!�B!���!�B!$�00"�B!�F�B!������B!�xB!�B#B!�BH�a`D!�B	<�!�B!���!�B!$�00"�B!�F�B!������B!�xB!�B#B!�BH�a`D!�B	<�!�B!���!�B!$�00"�B!�F�B!������B!�xB!�B#B!�BH�a` ���Yb3?}�&&�Y3�B�T���v�ii���}����{�7�HVͩ[�r���ַ��w��SN-����V��m�B�� ��Sd�d;���XL���[�� 0��MTƭLl䱗O	!$5�Y�"0+Aҩ6�!#B�#B!�BH�a`D!�B	<�!�B!���!�B!$�00"�B!�F�B!������B!�xB!�B#B!�BH�a`D!�B	<�!�B!���!�B!$�00"�B!�F�B!������B!�xB!�B#B!�BH�a`D!�BR����F�v�d����o``@V����?���rՌ2�-]��O<��=�7Ʉ�ܘ���.�����!�BHʑ���{ut����s�c�Zƃ-��VB��HO���tIKK�2�=����?�evV�d��!��W�����=��k�vy��}���|_����ѯ���O�l�ĭr�3�Zq�����v�df�ך�v�}�Z{����z���y��ׇ�`쯕BHr`` O�TF�Kldݼ"��S��W��#r�=�.�2��~�����T�m��;�s^A��"p��#\R�-U�2��@�ײ��Oj/���6ij��Ȝc��yYR��`Z��f_��7�u���&il�f��H�R�@��פ�<�[U��xg����V}��H_k~N�z�92gJ�L(��A�CK{�T�m���.iV�A�A�ϵ�8GM/�����	�ƅKr�\�4�Ϡ=��-^+��ά,�)�y:@rh�앚�r��]}=����E�Yz���,���˯g}K�Q�ϵ��GR��ƳJ��]l%s�=������_��礹�Nld��%J�W��^ӊ�l�<*�2!�D�6
!I��Q�HO�Q���\8Al�xi�����&v������'��n�'+�V���z��G��"
8���˟\7[��4K��o�Ǜ��;�?,�:����s*��̗k�T��L�|��#���3��>�@ ��kf�=�ϖ)*84��֓�'�	x���!И��w�a��a�T��]h��=uD�����覕Ur�se^U����sV��#�ډƈ�R�'��_?_��8sD��2h��ޓG�?S��	��b�~����)�����(��k;@j��BH��p͢I�{��Ie�iM��-�*]�U�W`��ˇ�Z"7,�rEEǍ��8W9��_��p�Y�_U"�~�J�:���sU���o^,*����5�U����<�c�������g���￻C�6�{�֡J���FfM.�'>�o[(�9���lWC��m�L�n](eE9�����):��ן�}������}���e��2Й�S���7̗��y���W+$!������B" /;S޸vZؠ�N>*5O^ҭu&n^5UR�a�"�s�U��
�L�Rr�3�E����}'��#�r�t����[<)lP�j�}�_m=a��B������w��Jy~�9�s���sW�,�ש�'\P���g{�B�g�A��i%�A�C�
$�^+�U��vV"!�\��!�D �%�,���,�Z����h�r�ˋ����0���X.7.��=�M,�yS�=��*��1)�`�a�U�����խ?Z?=�{V���s�=���\5�4����[!O�R�ݺf�nS�Tש���!��#B����� �0�4W��wu��([Ow���2 ##]ʣ<��oQ��}�P�H@%(t��HPw�X�fyU���?��)V��T�8/��iT����@!�~BH���]��I��M�Z�0�%M�0�%m��m�5�&Co!��00"��8��OB?}��Bb#B�q)�F�B� #B�q	T7��?�q)o�+�e�L!~��!�B!$�00"�B4��#�� ���B↟����~`��z	!$�00"��8ᷰ(��_!$�00"��� �!�F�/�4�l N���2L���Iw��vG!$�00"�B!�F�7��k�O;��D��?!��F��;b�h��y�W�!�� ���B|���:�{��ٷ��B�#BA��G1?K~�HGt�i�#;N��5��5K��{��C�s���g��km��m���w�Yu�sƟ����?;1��^lꔺ���������i��Eu�Ξ>�y�N�֓Ɵ���I�y������%��������3�z�[��"�go��:uI�֣Q�����!������BF���(^��_;��w>�볛cO�Z�'���j^+x�ӱ����>�������7q.#B���W�KFsu����]'�W_�*ͧ�c�Z���^�"G�sb�:��k�T��!�BI)^ٲY������/77Wdџ��w��G���b�Z&M��z[Կ���w�q������{{�E5��Ֆ-ٲ"wǉ_�K�����8�<��N.��yRl�8.w�\T,Y͒�b�E콓 ��{[l�y�"��K�)ߏ4X ��;;�߼��w���jjl�TY�l���^y	�   ���    ��   ���  p�Ą�'9$y���Z�"Q��� xBZJ��fkAY��R���w'2\q����^��Q��ّ`���ݽX_~l��3�XM���F�:Р��!+(��➙� L� �+�M�{n���W�hnq�r2c�3��K����V��kjIE�V��տ�pL͝� ��`��r3St��J}�%*�K��u�$'
����dݲ�T��{��7�n^ �� W3-D�ݱp�B�E��nI�~����B \�`��LW!sM�Y Ė�������� �J# �������4��.%)A ��� ���+�B  L�    �# ���
G ��k��J/8L�LD�`Hm�C ��`����B���O b���d]��{F 0� �Gt��W�N�i��B��9���H�6� `l# �V�ҧ�6W��0�I^�á�:{/o�	�s��;�?�x�P0�����Ы{��# ��F \m`(�74��'��o��+K���"������v�{/�8����?{i0�^r߀�̉��u�j�  6� W3�`���v�h���n�d&+)ars�S'`�D#�[ŷ� �#���PD͝�2Y�A  !   �=�    �#   1��   �Z�o~��m�Y���o���<�ߙ��ToK]��Oƿ-S���Rs��ۑQ�Ly+��   �Z��u\:�h���)�2S�a��[�  p�@������rR�	Gt��Wo;?�=  6��λ�3���ե�}M��d��}^��;�\����<��w���9����ZO8Q{ϐnXV�w��}�� ���z�zK+s�_?�V��;�*�q^k���Y��.11A�y��h���S��=��'[ �A��NeQ�>u�ݰ�x����݀�$'%h͂�qM���jS4ʉ( ���W�t�{h�<[FZ��f�4?M�� \�`���ӓ��,[ Ɨ���܌� ��`�#��Q%%�����B䐆�{�KN�k��V����_�z�O��OѴ��L0]��3�nN��̥w		�����zl������[�gّ��Q������G�Z�Z\�!'z��ԍ��[�T_���ɩ���Rh�o���ש�,_Nt�\��� xKj~���{�ʩ~��ޒ����w?�{_е�������Լ��v�*�l�����G�-#    �G0�Z�[l3��($ ��F \+dz=t� &��oX�mW�� ��`��z�u��[��!{8b ��n��[��V# ��$ ���FW�ڧ�w���7ϳG�p���=�v�^��  ��F \��}@O�U���4������d%%��n}�êj<?Zg`��#o.�w�w=��:p�]�5�pu��� b"p�p$j}����W�P�+J���2�u�w
�-�hT��Y�_h<����\~���H�PXC���t���� xB�f�LV�!�aY�f � ��!   �=�    �#   �=�    �#   �=�  ��P�d��F�I�͐�fp @l# ���������++=Y�Nvy��Q��0/�vc��̎+}�����ck'�3������o����M
��� b!p=3��-�J�ae��V�0'5��Gǹ��Oo�^����}b��<=�����c� `t# ������ז��[���YS������)���GN�w뙭g G �6�8S�sє�"���d��%zqG]� `#�/��K~p��[�|�uyݟ��>����h~i�V/����S4�8Sgz�zM���}��{j}���p����Gz|ҷ���k(�2`|I	�&'Nj^~�������k�!�SS&9�1  �F    @0 �.L�
 ��kE�Jo���	�
��7( ��F \k`(����m�
E5-}j�d��� ���pX�M�:^ۥ�sr�Jf?�}�U�� `l# �V�ҫg�T��[���T^�D�7�>;MP`���.\+Х޽�h8UW_P'��m�t�L�  c#p53'Ǧ=��u��J]��@Y���*j�W�Уg������#n����K�`u��[�����/ @l# �fF�j��/w��عN��Oz��G�̖hD�q��^  3�`�L�����,����'  �/#    �G0   �{#    �G0   �{#    �G0 �Ai��|ݸ�xR�	�"j�Бs��ke�E ��'d�'k��"]��H���.L���'���{��h@���zf��Y��Ѻ%���GVOj=�V02��<ޢWv�i�V��Q FG0�zJ���޿B7,+VFj���4z ����J�
2����d�4?]E9i��ѳ� ��`��L����t��
�&'N�:�����k�u�\��QZ� `4# �fΈ?r��)E��f�hie�
�S��=( ��F \+3-I˲���[0�k)�!�X�& �VJr��R`|��h"�D`L# �eJ� u  �#    �G0 ��F��� ��([i/#��^�-MS�7�5���,�������l}���jKZ /!p�P$��!
=`"�����1 �kJn��߻Ao��S�7���Ա�cr������q�ַx�J�x���`��z��:U�m���b#`L��}�u�E�C! FG0�Zf��ږ>m�[�{�� �h��+{�����  �F0�ju�}��g�^͜FI�\o`(�:+�k��r`�G����7���.�8֬]'Z� ����#Q�>٪/~k��}�\�9��Z��0�-a�D�Q��@���tY_�;#SRt��]*��g`X��A;h b#�sQ���=b/��~蜀Yce���A{ ��    �#   �=�    �#   �=�    �#   �=� O0��d�(/+E�ɉ�Zב�)j0;����s���z�a�j��o�ծ- �F0�z�IZ5?_W�蚅*�O}.�ѿ��ݨ�%�οhݢ�̚��$�Mn%Ѩ�/�[\�g���^>��� �����$�������Ԓ��)YgFZ� ���2+ݻ�R�M�zyW� �����)����^<e��+ -.��mkJ��:E"Q �D0�ZI�	�_��W��V8*�I���,U5� p%� �2�Ue
��L�:�� 0:� �2�^z*�  �<�    �# �Q�] �1� �VĪ�Ba*=`"�au� ��k�B��kP b�#j�P}[� ?Xs�M��#�������f��U��:e�;�ܫC[�)# �e��z����<�$K ��Dt��C�����r�r��70����r�{�ߞ�o��=ݦ�����`ϹaI�nY��ym���i�_�����Wȩ�����O��߬m��s���S�-QNF� /0�D�C병]E�#ՠ�O�m��S�����f �F0�'=�a�����X3?_Kʳ�D�[��L��꥝�Jt�R-��Qz*omp���m>�h�p4z(
����������Pu�vk�[U �Q= p5sf���O��~Zδk�';��)&��bZz^�Wo/NcN�ܱ�TN���z�N�uT�u�9ٿ�zJ ���'��]����P��N�'�\$�2�h�����k��D[����#   �=�    �#   �=�    �#   �=�  H�J��tNΤ�G�y�jZz��=$ @l# ��������j~����.�3���=?Q��v�fE�JF��-ӗ[;���ên�՛��ھz���V8 `t# �WQ���ݽX7./VAv�2R�[��0��mT)w��-��R��lN��g�˿�p�J ��� �ZQN��e���SNFʔ�3)1A�W��&���:Y߭�|BQ� `T# �6�$S�޶`�B�EE�iZ=?��O��� \�`��̙�e�v� ��$��� `# �������T_B @7Q ��`��L���  �d�    ��  0s�# ��`��L�7��z���5  ��F \�zU�LX	���s@�:��?, ��F�hT���g0�����G�:C�o�i1�i����Mڸ�T ���ԛ�io�  c#�s��O�޻�XN�s��W��g���huf����&�c���͚�^���3�_��ʢL^04Vs���&<���J���6�j�6m9Ԩ��> �F0�já��b��om�G�\�{��PA�½L����-j���sㅥ��o�t���_��S3�kEvP���S�d���mjֵ0���o}CN47�P��/��^���͛Bl# �g��U5��o~vP�|���ڨi_���bz����8R�G#�E�ϭ��h!����F <���p�Z&�����Q  ӂ`   ��F    |�`   ��F    |�`   ��F <!!PJr�R���8��R��`�$X/����G�^<���:QۥW���Pu�  �� �^rb�*�3u��Rݼ�D�E��ą��Ł���������_����%�k���M��D�zA��/-�s����[��I_1Q����� �Z���.*�]c�S!+#Y��%$�������F��ޯ���b>3�oF \mNQ�>y��)E��$Zi��<ݾ�L[5)����� ��9#>�4Sw����%'%�� ��fZ��' ��F \+3-I�J�`|��	�> � \��@�L\ �� 0*
    �G0   �{# �e� 6s� �P(���� ?���K��;]��GzN*�}Bn�X~���:�u�y�A��Ay��k�B��7( ���	���W��-�̽���hLWck��dQy���&����`��C:�У֮A�N�M��]ڴ�NLa c#p-S�ն��5z쎅�H�-�t7mh���oU���8� W�*���v�m��a��_Z����&'
p��������u`�G��@`��s�;�3��u�UoZ��tC�  �� ��|�}��!-*�VeQ��R&�v�h0[�k����� 0sF <�(�C��2Y�\���p�!  \��* �!   �=�    �#  \�k� �!  \�k� �!  \�#�oF   W����    �#�(�3  ��` �)X�{KRb����E��;'59��F"�p82���	k{�Vb8U$�Ʀ$%(�j#Q�ޱ�5������P8�pd�mM��5!�՚����V�o7�A��{\ ��` qZX��9řv��[��4�z_�Uiߴ��
G�q���kP�O��yya��T���v�lSG�И�_��PY�q]��7Ҷ#�c�_������ ���:U��?��+��(7-�pdr�k{�Ǽ?#5I�/+�;�=ծ��A ��` q�{]�>~�b�d���{��㗬`40�}&d}��k��2'�u���A_>�}���/)��Y�������ܬ]1��g޻\�����؟o��E����^�򂌸��k?ګ�ߪ��Go[����TZ��C�i���όy�	Z_����W�Ϧ��q��&��  G�5 ��F ���(�+L�z�e�{�nzl ��` q
hz
��N�=k���4�o�L 
 ^B0������n�Fnzl ��`   ��F 7][⪆=�  �!@�\6����i
\�z  �! �
�  �%# p����Mfz��� �=# ����v϶�  ��`   ��F �7���m�.< �%# �[T�*�]��ӳ��[ �l! ���5 ܨ�kP_������E���ǅr��٩�0%�D�(@��4D�N��. �=��^abF ���B���f�"1�7k�
ǵ�h4jmG��[����V���8�2`mk������=�H�~l���5�����aE��>_���'��m���x� 0sF ���>��)?;u¿s��;f00�a��v�^�?�u����/��4w���_���^oMs���B1�`u�n\Q��ĉ�����4�����ޠ����W�5�MU���3����.�]S��ԉ��tż�z|��tjIe΄��f�fzB 8����O|t�W��^~f��3������Z�7M��3�.U�����O����q�4�*::N1�G�u�tC�]�''%���C����vV�1iIx}��0W9�)�Ӵ>T7��Wc����#g;�b^��R�O1��^�[o�X6l�o�����_P&��~�Ͽ]��;��T�nX^��	���m�)+tƲ�D����
�)JL��2��'o���3&�n����ז++=y�u�V�CU�jh� ��F��ʥ��߸^N��7^�������jIy��h��*�ꤼ���O��SaN�V�Ϗ8:z���d������g�V����-�V?W%yc��@p��W���k�鶘��j�74h���/-Tf��E|wP�t�Uk[M�X,���)k[ٸ@�Ec�#�L�d����c�0�&-���[V�*7F@�ֱs]zuO���i5�j��so�����9JJ;���m+���b��]'Z��]��{]�
b���5-�f�f�n���B�խ���8����nN\���F0���U�w����h�TS�/i�3-@�:�͇�s+@t���	<���Q����÷̳[M.暡��~��v�6l�ж�>�j�p|��Z��@��	JdL�΀]��٭gu�yb�~�jh�cw,Pvz���\3d֋;k�˝�[�.8U�m?V�w�b;�\�����Uw����XM�����j�v�����
S.k�3�W�`��O�U5�u�X볷�z>�ZW���K�/�8kZ�N7X�l�9������(�ȹ'���޲>^����j�K���\N���b}�+ S�` WiϩV{)+�Pqn���-�M�^�����hL8zrs���Z��e9V�x�m�\���7�sM}q_���K���v+WYA�RG���7kZ���x�x�
<fYT����w[��jz�u��g��.Wkm�?���~��b�F��h�3���
M��C��0q�:�h/���0;U#3�	�'�P6�`�밂��~yB?~��d*sD����6-Df{t ��` ����o/SɌzw�n��j����v�a�0]`�Z�����\��yj��=?�?�� �"   �=�    �#   �=�    �#   �=�    �#   �=�    �#   �=�    �#   �=�    �#   �=�    �#����B�2���   f�h�&%hAI��eaI�R��$'���\X��߆#Q�#
E޽�5d}��1��-}��>����v�j��_{M^����&  ���i#�Lf�^��R/��V=w���oC��z���^U[�݅�܇�A0�&YiIZZ��Usr.�(�q�#!1���e�rߚy��|�;�w�N7��x}��5   ��ܢ��̱�5^Fjb\�HKN��Ѭ�i�W�>p1$���x]�z���G0�"�˲��4˾]i�!s;�L3aid`2a鄵����oiY \�Sֱ�ޯ�,?����V��r��[Z��Uss���<��`N��e㊢��3'�O���dûu&�`4	f'�uy��B5g�Ƅ�����傭�Z��Z�o��k  �.��m�U�ݺ��0�$�3���kK�kZ���xV}gz����d���w�ЍK
�6��ɛ:�$k9Z�-   ?3��L�dQi^��Ĝ���m��e�v��3'�M�!L�h��Ud�޵��Β��"�3;�������Nm>Ң�6  �O��\��*ֵ���ĽY>}��$���M���hk���ue���Ry�y#0�{�7���pD@  ^g��}����u�3Ŝ��
{�t�I/�kԡ�.al�1�_�o"s�/���˗�  �gy=�Ɯ�7��!dҞ��J�ˬ���d}�B��Ȁ���z���Q   n���ez���
D�3'�����6=��^�H� �����s��+����Zf_����Z�?�)   7�v~�>�a�+͚.��,���϶֨��\l#�oR}�
Ee.�d�\���]�z��Z5v
  ��L]�������`t�Aথ�z�
G\B��`�jN��Jd^�yc1��=��VOY	  �����Ȼ^Ix�� ���-������H��q�m0��-s���,�c�`~��E�~q���Z�N1�  p�%eY��Uߙk��P`��[��϶�ȏ|�L*6;�m+�3��t0o8_�d�����
  f��4��J�]y;��ch�37'��v���^9&�PĵDSü��;�+ ��f�Sߙ�t15Lͼ�<ۮ��:�"��M0����0�� ʬ���*�}  3��`15�����.�!�<�ROlͲk<?�E0��Wk�2X�N���X��xꨯ�,  ��q�5e���˄�e�ܜ�f�x^��`���Z���+�sf�/��  L3�g�[$�ӵ�<*χ#O�o����_�)�,�  �.��}�>q�|af�p��O&�+?: ��l0��nPa6c������m:�$  ��@(�]���;��A���.y�'�����6�$%���Xn�ӟn��X�  `���ana�~�G����E^�`d�(B�s����JOl# ��s�5��"�HI�d8�T02M{扂������zaO� 7����
�f��E λna����r�YL��nu�	F_��5v����\��`H�j����U��pK%�x�깹��'�
�djoS�{e@O#s����������X��0	,  �miy�Ut�������}������Ȅ"3| �/1!�Ͽo���'�U��'  �ј�V��W(9�����޵�j�	��W��\���^�"w)�M������!E�\�  .��w�ZaNa���8WM��zio��ʵ���k��Y��>��ۡ�_^9-  ��L�`j���޳X��W�)7re0ZV���޿Hp��Tiw�{y_�   �֕�5��t}��{��O|HM]�r�#3G�o߷HYi��t\Ɯ:�ܧ��=  ���"ۮ�ns�2�p�g?=$�q]�0;̚y���e�&Y��b}��  �SZr�]�� �w�������/��	W��n_Y��__!xǪ�9��m��}��b  ���LM �����:Rӭ�G[��	Ff��G70؂��u��V��K  ���"�ϣ.�x�;F"vM0z��9���C������G  ��� ���ء�z~��Fn��`TQ��q&��n_U�-�Z]��
  &�\&aj x���oU}������$�܌d�����
  ��I����M-��/���9>�_��ח���V  p��L�?L-��X��Tu�����Q���7Uj��&��  �� +�>��?LMO0������üQ>x]�~���  �7�c�9��?.��;N�ɩ���L���/׋{h5 ��L z/�I����	FW��"���  ȿ��j��`Dk���j ���Z'�92�ZZ�  �Z���V#G�;W3��{�)����"  �`�S��& /3E7-)P����ˋ���f  w3�tslL�oj��>g]2�`d��T�mfɭ+F  x�9����M����F9��ȍKi-»6Zo�s�2T��/  �N�X��`�L�O0��$7�nt�­ˋ���s  �d���H��7�sנ��Q��<@I�	F2g�~��` �[�Z�˙������S8*э�Y\������L�  ��\o�ͱ����	F��LMҚy�F��2�` ���K}�љ�FFJ���a9�c��5�s���(`4+��  ��jN|c�V(25�SN~;&�� �u�uF  ���Z5�����z9'�̊G�Q   �3=��1˵����g��F�l²�l�\3?�` ������@,�טSz9"��	�xLw:�.  �k��0k��iǩ���g��t��,-�VJR����  ���c��R�����X�`��&�<?]g[�  �����pJpD0�_�)`"���F  ��9f�,0����P��*`"8� �;p��D�,`2A�PhV�cփ��b��a�8� �;p�F<L&8R�=��0����Mgp�> ���	|��0q�} �8f#N������> ����#)%9A@<�Ӓ�38,  �L�X��	�`փQj��?p���$�  f��@<��	f�U��D0B|�7�  �"!^)#+&���t�� p2�ՈW*]�L:L�B �l�/'d�Yզ�b�8qA'  �Ʊ�J��H\c��q
  g�X�x�p��ED8B<zC  �ű�2�`���:�� ��q�F�F��ሲ�Lg�  p6�Ո���mփQ0���l p2�Ո�2����C�g�  p6�ՈW��tփ0L0B|� ��q�F��t���B#ć�P  8�j�k�#��c@k��
����!�#Q  �2�js�.�N0&̶YFU�}&��}P  ���1�`��rB&��`T�L0���;�l  �9f��O� LL5�H#ĥ��` �p�F<�	FRW���{�*�J0�d p�٘(�L&�m���	F��� ��1Q��A�`�~Q���4p�	3�;{� ��q��D�F8Z�-`<�{żW�	��  ��c�ilaI��X��8"9������  p��V�G0�x��8#8"u�LS��f	�A4  �bN~?tC�����Q�`HN��`d��&!��ut� �M���pP� �#s�g0��0�#  �����N6�hiy��ј#�pL0�b9Fk  �dNn�0'�rL0j�����9.w��9g  �ę^A��R��Y�3��S8&�Nu�p���!�>�.  �>�N����T#�:�!'qT0�y�M��s����k�@0,  �>�n���r��wG�S����Fk��
�`��f
  �k+��15�����Q���q��`���Ns���9  p3s,��7F25��8.�&�ߺw� ��"  ���	F��i����s���s�C���f�$o=N0 ��1���Z���D��L�oj~�q\02���<ܬ��!  �3�tsl�u傿9�G�#�ы{�fIy��_/�i  �sl'�۩�^��w"G#�%��|�R����ﴑJ  ��c�K{	G~��^��vl0����h- ��h5�/'��F�F�Dk  �E��9���pt0��ȟh- ��h5����F�������	��ܮzZ�  �8s�7���n�����N��`���Fm\Q�������o�
  x�9��j�x�Y)���<�n��N��`d<���`�OY�sc�  ���c�9���}�o3���"�?�Is�����S� �+��oz���#x���M-��Fͭ���vB  ~dj��<�J��]&�`Ds�w�q�Y[��
  ���L-pך�[�v��k��a�[�[����o0g��V#  �_��vA=�<dשv�]&�`d�۫g��>�V���8^`�Ϫ�>  �2���	����ն�;�<%�q]0:�ҧ�zZ��C+w���q�Y   �&�_����:Wp�p$j���N��4�`d�y���q>z�<���>٦�Q%  �Lm0�$C7/-�Ʉ��Ur#W#�oV[;N�6,c�q���A}��3  ���g�4/Mp�'���=r+�#��E�,H�ܢ�=��V�>   �˙��
��.[����7��ķ��QCǀ���c��'�*'=Yp>��047  ���
��	����	�w��W���I�����q��W������\'8�iZ}��\ ��r_��Ғ�[�.�k ��y渺��v�F�Ѻn���;�o|����Ex�����$  ��������*g�ƓGT�⍩W<���g;��~vX_��j�Y:�'�qP   ���/OiYE���Y�����sƝ#Ѝ�3���~�M�{�J���&W'��v  �j}�{{��W����W��M�O#�m5�-�h�մ��s��K   �����J?�ÛU��*̮���q��Pdx.&����.fǖc�v�S  ����[���ut��E���N�:O#�=������+1! ̜��ӿ�rZ   S�t����V��E��G����.y�g�����fu����[��\fO�	?�R��Q%  ���'��?�g	��͐ڶ��3�t��G^��`d�>ӡ?��a{���#����U驷��  L?3Z]S�~���F�O�뻛�t�#Cr���`d�������w.�Go�'L��u=���U:x�S   3Ŝ�=��k����뎦�O�:��Y-��E0��<�'��<����=���"��z  0����W��]߽�z��M������v�U~�`d�'�TC���ܹ�D�:]��v׹��7
  `6���z�U���]�r3������f;�t�o|��D��Ϗ�hm��8WE���75�C�W5{��)  ps����-su�N�ǣ�gHOl��/v�˯|�.0O����v8z��r!6$��^��>kV  �aN���3��9�0G+�������EM]��3_#ü ��œV@j��.���+\��7h"F�  naN��ћ��)?+E�ԡs]v/������E�a�_�v��4G���<�s�����;�}  ��9�k҇��ļG���̎Z=����#�.c^ �6�k����2���sbؗ�6��=:��+   73'xͼG��oԃ������y	ECǠ^��h_���.E0�y��t�9=���b@�_�!?   �2��?�pҮu��ζ�_D�C!at����;j�zL@���R-����af�K34#�  ����Lᒞ�(�9QߣW�7فh8b#M�y!=���^�/���E���1��w[���0яc�  ��~��9m\~��s�@\f�I����=U����d^`f��oV_܁�/ʗ[�Zh�;;ˡ�.  ��9A���:{Y37׮�n�����u��L���&!~��d^p/��q��t�[m�D+*�u͂<�;�%�LS��t�ȹ.�<�nw�  ��̉c�����/.�J��[e�yN���w0��Vmw��փ֭�6��!M�B�b\Q�c7î[����|k�����Yk'9�i��}�.  �x��om��(;U+��h݂��]�,�\|��;p��-��h��3a�Q�����t��� �����j���:�a�m��{m  `*��]��Ӓ�Z.mD��n���~�%v}���z��6�^���bz�f����Ŝ������wn�.~�e�C�[K�����#Q  `v��x�Y����0J��lߚ�L7�^S�ٷ�wn�9�=�F��:��    x�9������   ���    ��   ���    ��   ���    ��   ���    ��   ���    ��   ���    ��   ���    ��   ��`�f-�֒"    �!��Y�Zk)    ��	FǬ%�ZE�    2���Z��S�[�J    >b��	ki��Fk鷖
   �?�����ٿ/����    IEND�B`�PK
     ��/Z�I��5.  5.  /   images/ec55ee1b-9bfc-4adc-bb90-2198f3917cd5.png�PNG

   IHDR   c   J   ���k   	pHYs  �  ����e  
�iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 9.1-c002 79.b7c64ccf9, 2024/07/16-12:39:04        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmlns:stRef="http://ns.adobe.com/xap/1.0/sType/ResourceRef#" xmlns:tiff="http://ns.adobe.com/tiff/1.0/" xmlns:exif="http://ns.adobe.com/exif/1.0/" xmp:CreatorTool="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" xmp:CreateDate="2024-09-25T10:04:27-04:00" xmp:ModifyDate="2024-09-25T10:05:49-04:00" xmp:MetadataDate="2024-09-25T10:05:49-04:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0d4a73ee-b400-4bfb-840e-4582cd31f35a" xmpMM:DocumentID="adobe:docid:photoshop:102aa0f2-64fb-f64e-a33c-390250429f30" xmpMM:OriginalDocumentID="xmp.did:7c2c0979-bd24-4ddc-a181-e94452fe37de" tiff:Orientation="1" tiff:XResolution="1920000/10000" tiff:YResolution="1920000/10000" tiff:ResolutionUnit="2" exif:ColorSpace="65535" exif:PixelXDimension="838" exif:PixelYDimension="624"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7c2c0979-bd24-4ddc-a181-e94452fe37de" stEvt:when="2024-09-25T10:04:27-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d88baee0-672b-48c3-8fc7-826e592b23dd" stEvt:when="2024-09-25T10:05:48-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8569033a-e003-456e-822a-67d8550fecc5" stEvt:when="2024-09-25T10:05:49-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> <rdf:li stEvt:action="converted" stEvt:parameters="from document/vnd.adobe.cpsd+dcx to image/png"/> <rdf:li stEvt:action="derived" stEvt:parameters="converted from document/vnd.adobe.cpsd+dcx to image/png"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0d4a73ee-b400-4bfb-840e-4582cd31f35a" stEvt:when="2024-09-25T10:05:49-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> <xmpMM:DerivedFrom stRef:instanceID="xmp.iid:8569033a-e003-456e-822a-67d8550fecc5" stRef:documentID="xmp.did:7c2c0979-bd24-4ddc-a181-e94452fe37de" stRef:originalDocumentID="xmp.did:7c2c0979-bd24-4ddc-a181-e94452fe37de"/> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��9H  "�IDATx��|	|$e�����Nҹ�c2g�`.�`�E��U�p]�+����'?eWYWv��r\f�k���#s&�drM�N���������s5�����U��[�}�o�y�=?���=fdXO���v��f���FW�tw4��l�A�:V`Q5�	�4��xM�M�����cct:BcT%���I�3L�c��!<����(U���y^�ip��d�O����t���pT���qQM�ߩ �0��Ŏ0n�5�y�&"vt(�ؑ-B��(�_\8��
�$GE�7��Z�8<������3|XV�2Sp�;�7Zs���e�ֺ��q�f�1�bS�;z�D�Q�;���U�p�\vm�ַ8��McӒm��Z/���H0to�ec,B��B'�2'7�f�QE��Ǣ��j��'L���������(�m&��b]K:}֔�&F�<+��_@݂�P���>\>Ԅ�]m�с�I&�^U��}W:�[u14K6���ϫ������3;�`�B����x�fyL�9��ۉe���s06%��B^X����JC���l�P�A��=�g��ㅆ�I�fK��n������TVܸ�� ��яcC��xƅ��^�\� ��J9����7��;\FM"��ˊ��իL(�]E��B������2�W�r'18�^4��/-����p��� V5��ߋ�e�>MQ�	�M��G1�JD���� �;�����0vw��V�f�
la�}�	�Y�!b�����C�w{����0<!�0��{�,�,���:���(q�27�����`%w�h�[�kI�uW j- �h��k�*|���H#h��s�&���E.X�V������~'�ڄ�6�@�Q���4�K�]�X�:���)�ךed!�Mx�,��E�ɥ�ν
QK����	{ͥ�}���	����iq%�G/*����E��2��sp+�y�mZ�$���,�t@#�Т�������Z,)�ƶ�q+bR^V�1	B��qYY]���~K�o.+�X�����>%�K*�RcL�0�R�cNEb�|])���3r�k���0��B����A:?���ĕ+"�Ϧy�t�YE1X�K+L�\�;�0FI%���7am������EmE!b,�$.Qhv�K�0��m^?Yp��(����t㸄���"G�x(hIZ^J��$ii)�))Ϧ�GI1�Qp���ٌ?���)��F+�O�t�N��$a��p=����>1q-a�t1�nǡ>s���m{z�1�4��ɦ;K�f�X���H�Leְ�`��C܁��+�]�H'�)��)�`�����-h�Fьahl���<�� ���ϻrg����\EQa
�e�~��˷pfÉ�J�)(�uImWL*b����U�YY���݃XR�fv��B����D�ۖą�qd����v8sj&���	�;蚖M�&���Y�+݋����%��("�Mxc_'v����jɇ��=�/����W�B����(<���վ(��3�ط�E�ʅ�z9e+�"�NY{�b���dPK0�W�V�lG٬e4��B��K{��4<��o�����]���q 7Y	�at��yx������-�?�K�y��Uņ;���{��5�!㏪��A3�ߎ�ڥ����{����>rQ����d�w��q�nX9���%���t �>l�Sh�4��)J�� |�}?敨�c�ھݞ+�|�D���v�`���n���L�moRj{�?gR����ET<B�ʍ��)�mBYC�1�'��|��A��v 7��AB1���V[�r%g��;���������8T�E���!�~*.��ٖ����`q�1	�b�.�s*.{����op��m�ʳ`x,�wOr�횖1j�8������х,Im#x��)��Rۄ������~fc�L���%e1���;���F�&7�d}L ����^<��<Qd�T���2bÿ��a��UqeSA�<�����1�+@s�,&C\�!���T�FcR��å�mǑ��3�CUͩqQ���v{�!\4JX8�0��E�a�P�j~	�
��Ȧ�a4v�I��K#J�RY�ĵ�kP�2��탈F�+�ŕ5+0䥸�����u���]U��y��x��W,.Ñ�A��!)�k7k�U�CU11c���F�,�-@Ea6\�94���:�r��hN1��*Ʃ6�4��g`���lX1�N��w�4o(�e�l,���j��߇]2S���+�ER2�D㏴ྏ\��<�X{Pܟ�����^��O}�:���l�N�Q·�4V��P"�Vf���KuWݳ��D��,+6��MA3��϶a^U>��݊����m���i��J���U�d��#�DY�F�BQ2q3>pa^�Ԉ��C�	"�K�_���C�y��p4� �/�-���>���H+���Ɩ��6�*�Y��,��`�P�}d�-���GI!�b�F�&��$�u�����+�B�D#a��V�<f�CX@��K�"Q8+��C���]`	�,*�yac�5����������h&|vE.��#���fX3��9���;��D���h��#�A�� 	�dL�^]�����ڭ�m8��x�p��z�����������Q�8ō�|A\��䦘�Az�&%mjҺ��\��#(p���@R=8aþ�h��K�Qpj]C��zR��'�)%��a4��xukS�I,�����\P��l;eU�n-B�)N�4�����gI�3��!B���֟@��.�E��T��,��8�W�~}q:�S��	��%UB�^��������6TCa��ۏu*�3��H���lܺ�'F��ef��`�v�]�>�>���F��r8)Z�Z3�-t��X,)����hH����E�x,�<��T��\ ��'�	�jZByIA��С��R��zM��2�2��,j(Q��f�<{��j�{�����[SICYk�������i�!��!?ǆ��h�0�tH0f7U�����'��g��$��lg�^��+I���U
}s*�$����L)��=b��f����Gi-c�. Ϲ䦌��>����܁S��	c���HvS�AL@.e0�#�����t-瀹��b�R+�"�p���`:<���pUR����R$�'�W1Ć�L��W�r���p���ഝ��@��'��<��6�|~�1�L����HTJ#��QQ�YD��I�7��54��Jo�;�ԅٱ<�ֺ6X�WB���\r�ܭ�I5�dw)�3S{��(��{8��������n[VR(/�&k2N���r���[2���[�U����3��	��/�5�,^�rY�U{����}I��1�Y� ���g�8,g�8�.mf������<"�3�(f0�9�c�[���spl�uZq�ʙ�	�S�`2r;dE삗�,"���gD����#��S��H�˿B�nf��}��no����|��C���IƳ��0��K5[鎣]���q�:�-w{��1�:��	#�����>�l�=��g�� ++W��ങ0�j�	B��+R1i�`��V�"�_S�H�_��4m���~���8��(�3��[�t��dn;�9	��ȡ���3ـ�OPe��\����~2�pD�Z�;g ��(z�����F�,�A�ǔă�� ��"�]gKWTˈ@�I�k�~Y����,E�/�t���=����W͒kl��}r�{���-qI]��3�&v��?�3k�o`>ry���-ɖ���A�y_|z>�ژ��]wM������N����U%�i�kH{�
��2��?γY�E%#�6
r��][��dҋ&���h;�t���5b��m���o��$5
��	���X�Tv;�s	��V���d�u�we;�,�)yN֘�gܳ$.$�ȉ��V1�	wL�.UM4C5�ä�7�ɜ���4s�d6���qƄ��YT"Tˢ	�ċ9fBx����~S֐8�.�����F���e�6���F0��r�z��*�$���4v��Ṋt!7ۊ͇zp絳���A�ˆ�e9�ÞN|�4w?i1Å��ږ�������_>�\K8�r���f+����X�Fك�W��W�lAd�����vI�7��8��{���o�?��ى�}9>z�L�����_�u	���[qߏ�I�j!��y��n�� N`X����ֆ�,�Y
��_��P�%��Z�#$�;IK|��h��%��pוֹEC���Q�����~]3��s�w߸s±�XT��.�Ɖ.���xb�Q!�7/¶�h��$�����蕗_Cd�W6O��-ųa]�=r{����ڝ��C�W#���`t|��Ť�&Tg�8� �E#�H\m���ҐX.�J�qF��Jm��FE�#���;�"� Mv���q*�l�U4�q�j99e��%�ǉ�FrOF�:��r���6�ɂw�N�@w;:1���f|��p��q�t��\����D�O��f�V��Nl6+��r���T�UpUI���ݤ����e&��X���S)�9��A������19�x�����:��3�E^-.t�~�+���_$yZ%N��$A�%�^Pr�e��&iS�1�<����&i�3�����~,��ݸ����;����E3��B�@�w��=<�;	�ld]���~���a��尕�,ǿ~�0"�
��ƔA�OFlʜ�>򹕘[Q�j����Ō�\���qý?<}���?W�/ģ�\���>���h�f��5QLA��(*�Zj&�{1����J�~�c5�����k*�N�݂
&�_-�L��l� �H<[r�Ŀ�1�@$��������{6�"S��`7>��w�2N�IJ%�GF����2E�{�2=���EW�㔍�'�ɎE(�GB;b�7��9���h��� T:V�����M'�W�,�'���-g-O999(���}�r���0��s�c�T�&�J�m���W.)������a32���E�⛿؋��0�����E�D$�n-����I�s��X�BO1�$��7�Ɓ�l��c'�v�-��t"�wLZ|/1�#y�M,ڂ�H	
�	n"��0����	ސmRq�{�B�n���+�4����g�Q�热�b��Ћ>^�����d��|v�f䡄�9��b��RU�[T��u�L�kq㾟���_�{o����
���8��f7̮:�jg"���'�W�h�0�Q������w�rP�w���T��9[��2L�x��H�씥����&H�ZS�p2Q��Zx�vL�9U�S=�� ��P���V�َL��V7~��!x�M�=AQ��l'r]9Iad9��;gY|��&�b�IfE�o6�d=�EtR�0ީ��.?��3�8#��������m}>8mf�~W����O�p@�{r}��tR7{�rL2#��x�j,���c�zx�����/]��o���^���z8�j�9
�cay���n4uyRӵ�{���8i�	d��yNm*n���&7��r=�D��k|_éL��Z��������)��{����-l;ҋ~�Uj��U��?���t�t�l������M�iz�鮥�{ŷ��;PY���Lo����J�=�o"�����KZ�zݢ��K]��m�e����ßL�!o�Rfu��j,�W��]x!CSs�j����ei5��z~��Q23,�6�-����ɷ���À��-��'��42�H�)|��;QT�BÖ��ͽ���/=�^�(z���.fӭ��ȯ��h�ZQ-�s��W����6J����X�,�M��E�Ξ�q�݂�1�&i&�[Ϊ8�s ���.�x�у8�>3�\��O~�:�<���w��㕸51H�{hu7�J1G^�K��΍F�j�͎0e^���94SL��t�&��Tȸ0��7������&n�?�F#|�0�ᖅp9-��4���v�@�6|�f������6e'��� ��^P�Ì�fI����f:��=+�/�V����w�p%�����E�x�`?�񹣓b�^���=�إ_ǁ�#����)w�g\luU����W�~��E��YZ!{xy������j��gf9�c�=4S�.���h�dmīv��r������؏������o��eY}�ʄ7�wa��>X��B+//E~���1G�]/..BA�lT�z��!d���
�ÉA7�54S��/��q(�ܽ=0�,�aB}�!_���ߑ�p��vl��g3�W�w];}C������1���Xc���+�I����twK8��A��2
<� y�Q��L�Lu_�a�ˍ�?R�f�ᵗ_�ˏm��D_ψ,��,v��������g�
��TCU�
J��bA_��m�B?��D�pz�`7���	�]�r�~��g#<�(���}t�>�S9��ձ����
�kY�;�H.�����~�O���'�L�t��k������n��L�8/~Q�����x?!S������p�KQ��Q��3A�_�c��-ÿ����̠t���WQj���}}�Q���E��E��h�ҽ�k�Z�E} }����� ^8t90�#��Q���4k)�Oj�XS�+az6��I��즥�3Y�є)褪��ݝ��ϗxU!�_b���ƞ�����+p2R�c�Ͼr5r,�^�� ����
��B|�?6c�`���O��Љz��zY3�6Rf����*٘�*�&�rΤ��HfF�������}�C!�m��+On��*[�Ú�-A�����pGG�d��	�D�V1����3Kv���0�3��U�\?
g�%��nÝ���O���-���a�i���-��~���~��Puk+��Ex��}�~E��T~����>��a����LUM|"�}%��8al��X8Kx��\�|6E�x�,H�5T�r��k��c3i���)7K�'J�s���\|�,��[���W]���,̛Q,nǕ3�9U��=��UE�*�BVv;�j�Q��As�NG4��'�����`��e��eR�s�D3���9�ls ���~���tɚ}�6��x���H2.Na���j\��)�յ��������t�z���J���ut����n�������6���ۋ������v{�v[��.�]#xiK;�xsO��o~���=�:4�]>n�[��Qh�:���zB�'��tm1�&�:��LYߠ��2#��_ ���� �
\��h�%W�U	�j������o�&aҩ^�'�X�h!n�q��y�ť�4���'���eO/�T4YIs7���/M Fx'Z[����^:$sqb�էwɹ�^?��8���wJ���w<*��8�L�+p�/@v�+��d�W��x68
!;ϑ��z������wX��+w�9S|��*�wV�
���;�\N3*ySV�M&v�B���F�Do)|�h���x��R�u��#����z;DӃ.�C��TY	���YCǟ1��-~n����ÎG^�T4]S	���Q}��uj�K��������-YD��N��*�
�϶�0�F�854�XD�|���Payي[.���KJQ����:���0v4��8�7*m�طt�)�C�F��^9<�|bQ��^�ן۟d�����4F	�W~�g��h����efI>����"/���{��a?ީ��ZJ$؝����	V�����1�\_'f)'6�2$�_\�+�7���ޮd�3����$�O �GU�7	�������l��gz�7�;<���T`^�|Q>����'��wDjr���oM�Kׯ����v�:=)�0M<��J�����RT����&�"�n���ԉ���ӕ���pT��5���}���$�)��N.����N,����?���D`��yE�|s�s214M�D���*���w,�?>W�F�mS�m�7
5b�E�˂HH7�P�
>��9h��r�n���6w@��Z�k.�9�6O!�5-����)�[W���n�#ǩ>�2��E.���|������/'	����+��2RI�~���g�ۿ=�L $H�F�Oz�~�ߧ�Lw�,x�Y@���r�v[%)�!/�XL�fq�Iy*p��xN��?�b��{z,`�0�Lo��G�������ݧ$NGR��(c�.t��0���s˳��?�g-.�N�7t��`a����5(�I����aS�Zv:`�W�k������>��t�߮	�9#�D�a0db/V�ޑ���Ԉ|�|�_u��,f����c"$���*D�l,�����?�o�?`AtP����p�|^]V+	��]*_��(���~T,���kΤ��)�)>���~I�bѳ{�9J�kS����[:�bc�|(���� |,�L����j]����g���N)>���t��]��esE����(x�����kr&�I`���'�qق�x�~��=�MG��߀��&�Z��7P\]�<��7�練����ͤ�t2��Ηjg�ؒN��
�-S�v����4�����|��Ų����=��N�3hE}�������2�ޟ�{R�p~W�t�{���?�}��y*����x��f7�E��?�\���ާ�R{$��F��;��i�E��D���vH@���j%]�.�T�p�`��x��k�����������}?݇O�����Q�cMf~��$�����lm����d��/	d��x���mb%�_V���y��+�7�MG����v�����p=C_T	��u���0�,�yvy8�X�=n{��;�R������7_8��B'f�f��ڤ��;��Sa�]:^�]�K�Kp>��,%��e��_B�>H�hVPδ&��|!$����Op�ā�j���	�[XK,���TB����    IEND�B`�PK
     ��/Z�J�?& ?& /   images/fae5eb44-bbe2-4b21-a13f-fb7a66868d1d.png�PNG

   IHDR  �  �   u�c   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���=o\e����5c+��$)��)�R���D���
Ж�@84�l::`��d[2�5cd�E$,Pb@�tk�Z�����8�il�u���9�����5��+�j�֪~��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��J �����s|||�t    ��?��O����ڥ;    �4����� ��K� Of�t �8���{�?��?�{���o�[    ��N    �S�s�߃��DĿ�n�L�t @iu]��s��t         �/�ܭ������1pfZ�47RJ�?Z         L��~��j����3����JDlF���-         ��������!��1pf����ţ����x�t         '��h4��a0�܁��4������        �t�2�6WVVΗ��;0Sr�)"��Z�         NՍ������\����3e��x�t         �/��F��Y)�<<w`f�u};��E�         ��UU}T:x8��L�/���#"�n        ��}UU�ۥ#�?f�L�����V�~D�+�        @)"����/��1w`�5M��F[�t�         �Z�9������~��;0���Y���q�t         c�R���^�w�t��܁����ю�{�B�         �ʳ�v�窪K� ���JKKKw#�V�         �O��fD|��vmia�x)���4��9�Kw         0���t:_�� ���;0U�~3"��         `"|ZU�Ua��Sc8>�R�.|�         xxwWWWo�� ��(0�~��j���[         �(�ҽ^�w�t`�L����K)�_#�r�         &�b��z���v�t�:w`�moo/���͈�V�        ���9>>�Z__�t�2w`b�Ӆ�"��-         L�뇇�����ϕ�Ye�L��i�D�;�;         �9�W�sΩt�"w`"���R��t         �'�|{0|V�f��;0q�~=��u�         �Wι[Uջ�;`���i�)����+�        �TK1������Yb�L����+��K�         0�s�?��J���0p&����ţ����x�t         3��h4��kp܁��4������         %\�F�+++�K���3p�Z�9ED?"^+�        �L�1??�}�۝+���k����G�{�;          ��F��Y)����[u]��9Q�         ��UU}T:���;0�����)���H�[         �o|UU�ۥ#`�cg�z�պ�J�         �oH�M���tLw`�4M��F[�t�         �r�?���k�C`��c�i�ň�WK�         �C��s����].���툸/�n        �G�l��������!0܁����t7"n��         �G�s��v�]�\xB^"���i>�9X�         ��[�N���0�܁��~3"��         ��iUU.|�'`�3�O)}�E         L������JG��2*�����V��KD,�n        ��N)���z7K��$2p����үq�t         ���V��`mm�j��4������^h�ۛq�t         ����������S�C`��g&�.\��/�n        �3p���������!0)܁3�4͝�x�t         ����+�9�T�&��;p&����O)}R�         �Z���`0��tLw���u�z����         PJι[Uջ�;`����i�)����+�         �����WK��83pN������،��[         `��ϕ�qe�������GGG[�L�         #G���`0����`����i����~�'�         ��]�F�+++�K���1pNT�9ED?"^+�         c�������nw�t�w�D�����         �q�s~��鬔�qb�����o眿(�         䃪�>*���8�����zD��-         0a������0܁'�����jݏ�s�[         `������X:J3p�H�4��h�O�n        �	��s����_+%���i�ň�WK�         ���s����].���ecc��"��-         0E�m��?WU�X:J0p����݈�U�         �M��fD|��vm}�9z��5M�q����         0���t:_����f�<���ߌ�;�;         `|ZU�i�)��C�ϧ���         8+wWWWo����b�
<����m�Z�D�b�         �!�ҽ^�w�t�w����^J)��K�         �Zl�Z��֮���f��C����v{3"��n        ��9>>�Z__�t�&w�w�Ӆ�"��-         @\?<<����|�t�w�w5Ms'"�)�         ����+�9�T�N��;�����O)}R�         �k9�ۃ���p܁�S���9�Kw          �-�ܭ����p�܁��4͍��FD̕n         ~W��A���t�$w��988��q�t         ���s�?��J��I1p""bgg�����VD<S�         xhG���`0��c*��4������         L�+��hsee�|�xR�0�r�)"��Z�         �ݘ������Ε�'a�3n��x�t         �dr�ot:����$�a��u};��E�         ��|PU�G�#�q�Ì�/���#"�n         N�WUU�]:��;̠����V�~D�+�         ������K���2p��4Mg4mE�ӥ[         �S��s����_+���fH�4�q?"��n         Nݥ��^�r�xX�0#666�q/"^(�         ��g����UU-���a�3bii�nD�*�         ����͈�����3�<�0���8��a�         ���:�Η�#���Ô���͈�S�         (�Ӫ�\��X3p�)6�O)}�u         �?�]]]�U:~��+L����m�Z�D�b�         `l�SJ�z����!�[�a
���^J)��K�          cg��j=X[[�Z:���;L����v���J�          c�s||�����T��K�0Er��k�R�         `�]?<<����|�t�_�0E�����          &C��������s*��05����O)}R�         �,9�ۃ���a�S����s�_��          &Sι[Uջ�;��&\�47RJ1W�         �X)"�~���!�6w�`W"b3"Ηn         &�|����`�\�f��;L�����GGG[�L�         `j\�F[���>�"�a5M3?77�CD8!         ��+��hsee�|�f��;L��s��~D�V�         �Z7����v�s�C�-�0a���?���Jw          �-��F��Y)��l1p�	R�����;         ���AUU��`v�Ä�/���#"�n         f�WUU�]:��`�`�z�պ�J�          3'E�7�~���!L?ws���ϣ�h+"�.�         ̬���O�~�Z����;���i[�փ��Z�         �y�r�[�^�r����;�����vD܋�J�          ���v��sUU��C�N�0�����Fĭ�          )�|3"��v��Ȝ8���i>�9X�         �w���t�,��1p�1S���q�t         ����*�r��a����SJ߅w         �wWWWo��`z�����V��KD,�n         xH�ҽ^�w�t�������үq�t         �#Zl�Z��֮�a��Ca����v{3"��n         xL��������J�0�ܡ��s�p��ZD�T�         �	]?<<����|�t���
j��ND�S�         �$�_YXXX�9��-L&w(doo����'�;          NR���`0��t���
������ץ;          NCι[Uջ�;�<�pƚ���Rڈ���-          �$EĠ��Z:��b�g����JDlF���-          �l>���`0x�t��������ţ����x�t         ��8�����$���@�4�sss?D�H         ���2�6WVVΗa���)�9���G�k�[          
�1??�}�۝+�x3p�S����yD�W�         �����Ng�t���NQ]׷s�_��          TU�Q�Ɨ�;���p�rJi="R�         �1�UUUo��`<��)��߿�j��GĹ�-          c&E�7�~���!�w8a���ϣ�h+"�.�         0�r�?���k�C/�p���Yl�Z"�j�         �1w)����.�a|��	���hGĽ�x�t         ��Xj��?WU�X:��`�'dii�nD�*�         0Ir�7#��n�kی�;���i>�9X�         `B���t�,Ay����~3"��          �p�VU���g�O`8>�R�.�K          '�������c�����g[��/�X�         `J�SJ�z����!�a��aww�RJ�׈�\�         `�,�Z�kkkWK�p���moo/���͈�V�         `Ju������ן*��2p�G�sN.\X���J�          L�뇇�����ϕ����#h��ND�S�         `�_YXXX�9��-�wxH{{{倫>)�         0Krη��g�;8���~=��u�         �Y�s�VU�n�N��;���in��6"b�t         ��J1������t��?pppp%"6#�|�         �7�s�q0<W:��c��cgg�����VD<S�         ����8����}�2p���4������         �x�2�6WVVΗ������9���G�k�[          �M7����v�s�C8Y��7���?���Jw          ��r�ot:����,w�u]��9Q�         ���AUU�������/���#"�n         �}UU�ۥ#8�����[����8W�         �G�"�~��b����;3o8�y4mE�ӥ[          x,9������!<wfZ�4��V�AD\-�         ���s���z�K���ܙY툸/�n         �D,��ퟫ�Z,��1pgf---ݍ�[�;          899��m�۵��@�h̤�i>�9X�         �S�V����t�����S���q�t          ��Ӫ�\�<aܙ)������w��         �wWWWo�����23�~��j���[          8�ҽ^�w�t�������{)��kD\.�         ��Zl�Z��֮���3�������fD\+�         @��������J����3�r��k�R�          ��~xxxyy�\�~��;S�i�;�N�          ��9������sN�[�m�L�����SJ���          `|�o��Jw��ܙJu]��s��t          �'�ܭ�����=w�N�47RJ1W�         ���"b���_-�_3pg�\��͈8_�         ��6�s�q0<W:���������s���h+"�)�         �D�8������0pg*4M3?77�CD8A         ���2�6WVVΗ���)�sNя��J�          0�n�����v�J��:w&������^�          &W���N��R�c��3�꺾�s��t          Sც�>*1�ܙX�����zD��-          L����z�tĬ2pg"���_o�Z�#�\�          �J��o�����Cf��;g8�y4mE�ӥ[          �J9������!������4�b��zWK�          0�.圷z����!��������ю�{�B�          f�R��������!��������t7"n��          `v�oFķ�n������M�|�s��t          3�N��e�Y`��ث��͈�S�         ���iUU�R:b��3ֆ���)��³
         @y����z�t�43fl�u�l���%"K�          @D�SJ�z����!��������{)��kD\.�          a��j=X[[�Z:d�3v������fD\+�          ��s||�����T�ic��X�9�.�E�K�[          ��~xxxyy�\�ib��Xi��ND�S�          �H��������s*�2-�{{{倫>)�          +�|{0|V�cZ�3�~=��u�          xT9�nUU����4͍��FD̕n         �ǐ"b���_-2��)����JDlF���-          ��s�?��J�L2w���ٹxtt�ϔn         �pq4m���d�NM������N�          0M��F�͕���C&��;g.�"���n         �Spc~~��n�;W:d��s����?���Jw          �i�9���tVJwLw�T]׷s�_��          �3�AUU���$�p�rJi="R�          8#_UU�v�Ia�Ι��߿�j��GĹ�-          p�RD|���_,2	�9u���ϣ�h+"�.�          ,�����J��;wNU�4��V�AD\-�          ]�9o�z�˥Cƙ�;�fcc��"��-          0�����UU-�W����q�t          ����͈�����r�?
��i��s���          �1�V����t�82p���u�fD�)�          c�Ӫ���tĸ1p�D���SJ߅g          ��1    IDAT�ȿ����*1N��91u]?�j�~����-          0�)�{�^�f�qa�Ή��ݽ�R�5".�n         �	��j����]-2�yb����v{3"��n         �	�9>>�Z__�tHi�<��s�p��ZD�T�          &����������J��d��i��ND�S�          &]��������s*�R��;�moo����'�;          `Z�o��Jw�b��c������ץ;          `�䜻UU�[��wY�47RJ1W�          �P��A���t�Y3p�\��͈8_�          ��|����`�\鐳d��C��ٹxtt�ϔn         �pq4m������P�������!"f�          ve4m����/r��C9���x�t          ̠�������&6����f�D1� ��酁����"@�Y�@�E��⦋$��.���5�vm�M�U(�p*���P��-pqa�c��EQ�%K���2�9g^�y�$~��g^>�%5s�+�Cj�;�:th.w�n3p�}-//7"���          fUJ�Kx2w�n3p�=---}5���;          �xbaa�OrG�&w������������          DD�_/,,|-w�n1p�-//?�l6��          ��w�ȑ����������������-          �oؗR��#G�|"w�N3p�W��퇚���X�          �]=�Rz���Ï��I��رc��x&">��          x_[��O��S�y����_��          ܝ��g"��:4���K�����wRJ���          ܳ?<p��_��	�����W"�{�;          ���g�;wă2p�q����n4��          `�����/�xF�3lii���f�_#��-          �k5�g>���!���}F��⋏4��Fģ�[          ��P��|����z,w��0p�AǏ��j����O�n          v܁�����?�;�^�Ϙ�Rc���OE��r�           ����p�����r/�gL���^D|=w          ��RJ��o߾�SJ��-w��}����K�l4��          �)��=z��sw�-�����Ŕ����           �VJ��������3��n��h����-          ��kD��#G��A��c�>�^~��E�s�p�           ����?=z���Cދ��{�><�������          d�Ắ�?z����ܧT�ݞ����QD��          ���X]��=���y'�S(�Ԉ�#��-          �������?:th.wȯ3p�B���ߍ�o��           �SJ�Kx2wǯ3p�2KKK_M)�E�          `�=����'�#���}�,..~��h<��-          �D�녅���x����X^^~��l�8">��          �����#G��n�������Ѻ�������          L�})�9r��'r��O�v��P��|6"��          L�GRJ�>|�ќ��رc��x&">��          �x[��O�`�>�<����r�          `:��>�С,[s�	�n���R�v�          `����2��O�����D��rw           S����^�����Y\\�t�����o          쮿����|A#�	�����f����P�          `���3���^�����x��i4?��Gs�           3�f���SO=��^����8~���V��\D|"w          0sTU���O?���~!�1�Rj�߿����\�          `f=>|�ر�����v�����z�          `���~�ƍO�����c쥗^�f�����           ����G���n]��}L---}1����;           �.�thaa�v���c��n��h����-           ��G�9�;}a�1���/,"����s�           �����?=z��;yQ�1��/|x4=���          �}|����=�c�g�1�n�����~;z          �.�X]��=�������@J�G"��[           �ѧ�����СCsz!�1����݈�F�          ���R�ҁ�|���g����Ք�_��           x@O,,,�Ƀ\��=�����7��#���          `��������Ɇՙ,//?^��������l;}�����o�;         �7�f��v�ڇrw o)���?����^�h������G����X�`���V���W����E        �	��}(���rg w\k4���O���'5w��w�n�j6�φq;���,���q;        ��*�"�Ν��HJ��Ç?z/O2p�CǎkE�3���-���p+++1r�         ��z���;����V�'��������_��l��:VWW����N        `���(�H)�N~)������C���v��}����樂����c}}=677sg         ���6r����˻y`c�K�XZZ�J����pC��W^y%^{��         ����طo_��W}�[��֓�� �]�����f��"��-���/���z�         v�?����>�;��J)��?��?~���D�]�����f���a�c����q�ԩ�         �~���(wpG��h<s���ϼ��wɋ/��H���iD<���v���8q�D��r�         �G��0r���P��|����z����}?~|_��z.">������cee�R         fPQQ�u���UU=���O�����}������*">���VUUt:�����S         Ȥ��EJ)wp������ǎ��ۿh������"��;�m)��v�q�֭�)         d�R��(rg o�R��7n<�Rj���VΠi��K/}3"�*wp���z\�z5w         c �UU���|�������\��'?�ψ���=�������F��/1����ꫯƫ���;        �13??���˝ܑ"�}�[����n�?��n�]�|9N�8�;        �1�o�>'��x6�/�?��_~�c��腈���-�����XYY���s�         0�>�����\����V�I��/|8"�="~'w�������JTU�;        �1WUU�Z�h6��S�m���S�ݞ����QD|2w�m0���J���)         L��REu]�N~���>��q$"����V�ut��(�2w
         �͑{J)w
��eyy�����'N��7�x#w         �����zF�0Z�&����W#����l��؈K�.��         `�����똟�ϝ3���,..~��l�("�r� �^{�8{�l�         �@]�17g*
��ߥ����#��"���-��+W�ĩS�rg         0E���f����-���w?�#⣹[�m[[[��vߺ[         v�h4�V��f3w
����n�j6��F�c�[�meYF�Ӊ��r�         0�ʲt+d`���;֊�g"⳹[�m��0VVVb0�N        `��������3p�~D|9w�����v����r�         0RJQE��r���0p�v�;)�o�� �X__��7o��         `��um�{��;`---}��h,DD#w�����q��         ̠�R��bnn.w
L=�_�����f��\D| w��q����         ̰��#"��a�������Ǜ��D�Gr� ۮ_�kkk�3          ���f���	.�f�q��/>�h4~��n�mmm���j��r�         @DD�e��(wL-��8~���V��\D|"w����G�ۍ��r�         ��(�¾v���SJ����?���l��*:�N����)         �������sg�ԙ��{���^D|=w�-��n7nݺ�;         �UJ)ʲ̝S��; ��^z��W�;�;�����ի�3         �}��������ϝScf�KKK_������x��W����3         ஥�""bnn.s	L������O5��#b_�`��˗ccc#w         ܳ����hD�5��\�Q3wz��/����x."��l�y�f�<y2w         ܷ~���0wL���M�^�pD�{D�N�`��۷cee%��ʝ         ���h�Z�l��԰cf���n�����~���l��tܱ        �TH)EQQ�u��X31pO)5"�HD|!w�����v�Q�e�         �1)���z�Rʝi&����ߍ�o�� �X[[�7�x#w         �8#w����mii��h�n�mllĥK�rg         ��I)E]�1??�;&�T�?�l6s�[�m�Ν�s����         �]W�uDD�͙��ݚځ������o�p�`ە+Wbcc#w         왪���hD�5��]�QS�NY\\�hD����n�mmmE��}�n4         �UUE�Պf��;��ԽK���C�f�وx,w��,��t:QUU�         Ȣ,K;:�S5p?v�X+"�����n������~�� w
         d�R��(����)0֦j�~����Gėsw �꺎n�EQ�N        ������r��ؚ��{���NJ�۹;�;�����͛�3         `l�u��Xx��;aii�+�Fc!"�[�m���J\�p!w         ���R�u���S`�L��}qq���f��@�`ۅ�̙3�3         `l�u�F#Z������w����Ǜ��D�Gr� ۮ_�kkk�3         `�UU�f��ަ�;�~��⋏4��Fģ�[�m[[[���)��)         0ʲ���rg�ؘȁ������Z��"��[�m�~?�ݮ_�         p�z�������SJ����?���l��*:�N����)         0������sg@v7po��ߋ���� ������ƭ[�r�         ��J)EY��3 �V�{��K/}3"�*wp���z\�z5w         L��R�u���S ���/--}1"�1&��y�V���j�?>w         L���#"bnn.s	�1�v���F��|D���l�|�rlll��         ��SUU4�h�&b�;j���{��8��n�mnn���j��r�         �T��*�ͦ�;3��;���Z�ߏ��;�m�oߎn���G�          ����GUU�3`O����� :�N�F��)         0�RJQ�Ci�)��]��*:�N�e�;         fFJ)z�^��r���0p����Zlmm��         ����I�F��w�}mll�իWsg         �̪�*ʲ̝���xO���Z����3         `�F�����3`W���ʕ+q����         �/���3`���hkk+N�<)��)         �۔e��(w�
w�7E�N'��ʝ         ���,���J��������� w
         �.RJQE�u�;v��;𖺮���DQ�S         �����=��;v��;����x�7rg          w��k�2U܁������.]ʝ         ܣ���,���#܁�p�B�?>w         p���a�������a�]�~=666rg          h0�p8̝��f���V���FJ)w
         �ʲ���rg�}3p�U�et:��         `��z=�@&��;̠������`0ȝ         삢(����p��aƤ������۷s�          �$�EQ�΀{f�3��ɓq�ƍ�         �.���ȝ�c�3�̙3q�ҥ�         ��FQ�e��k�0#.^�gϞ͝         ��p�� w�w��������;         Ȥ���p8̝������۷���F]׹S         ����~TU�;ޓ�;L��`�N'F�Q�          ��RE��\ƚ�;L���bee%ʲ̝         ��7G�)��)���aJ�8q"nݺ�;         3u]�3��a
mllĵk�rg          c���(�2w�w�2�Ν��_=w         0�F�Q�����+�a�\�r%Μ9�;         ��� ��a�x��;L��7o���Z��r�          �,��F�3 "�a*E�n7�Ν         L��(����`��n8F����          �)��a�dg�����t:���r�          .�EQDJ)w
3��&TJ)����7�ȝ         L����(���0w�P���J\�r%w         0e����,sg0��a]�x1Ο?�;         �R��0��~�f��;L�k׮���z�         `����3�1�0A����ĉ�3         �Q�e�F���w�eYF�Ӊ��r�          3�,˨�:w3��&@UU��tb0�N         fLJ)����R�f��;���Rt�ݸ}�v�         `F�u�^�ȝ]g�c��ɓq�ƍ�         ����:��ȝ��3p�1v�̙�t�R�         �����*ʲ̝�3p�1��_�"Ξ=�;         �W���3�R�0�677�ԩS�3          �Q�ߏ�h�;�)d�c���E�ۍ��s�          ���,����Lw#�~?VVV��         ���RE�P_v��;�������DY��S          �ʛ#��R����;������u�V�         �{R�u�z=#wv��;������z�j�         ��R�u�e�;�)`���={6^���          d4E��ϝ��3p��._����j�         �1b0��`��C&���q���H)�N         �1�~?��a�&��;dPE���F]׹S          v\Y�QUU�&��;��p�NǝI         �T+��a��3w�Cu]G�ۍ^��;         `W���(�H)�Na���I)���Zܼy3w
         ����:��ȝ�1p�=r���r�J�         �=UU��;w����ŋ��^˝         ��h4�~��;�	`���ڵk����;          ��`��0wc��v���V�8q"w         �X(�2F�Q�Ƙ�;쒲,cee%��ʝ         06ʲ���sg0��a�F��t:>F         �פ��(�H)�Na��K)���jܾ};w
         �X��:z���;���v�ɓ'�ƍ�3          �Z]�QE�ƌ�;�3g�ĥK�rg          L����,���w�!���/��ٳ�3          &�p8�~��;�1a�;`ss3N�:�;         `"���3���z�^Y�0    IDATt�ݨ�:w
         �����1�rg���;<�~�?����0         x@)�(�ҡ�3���SUU��t����N         �
)�(�"RJ�S�������Zܺu+w         �T��:z�����2p��p�ԩ�z�j�         ��T�u�e�;����={6.\��;         `��F�����3�c�p._�gΜɝ         0�A���!w�K���q����          3����p8̝�1p��PE���F]׹S          fNY�QUU����;���p+++��         Ȩ(
�� wxu]G�ۍ�(r�          ̴�RE)��)�"wx)�X[[��7o�N          �/.�2w�����+��W�\ɝ         �یF�(�"w����������3          x��(��~�v��;��k׮ũS�rg          ��A����0wx����8q�D�          �BY�1�rg����ʲ������*w
          w�,K��)b�1�bee��T          L��R�e)��)� wf^]ױ���^/w
          ������zF�S�������7n�ȝ         ���:��0r�p�̴3g�ĥK�rg          ����~��;�`��̺x�b�={6w          ;h8�`0ȝ�}2pg&]�~=N�:�;         �]���c8���>�3sn߾'N���R�          vI�ߏ��rgp�ܙ)�~?VVVb4�N         `���(���:w
�����QUUt:�����S          �o��SJ�S�K�̄�R���ƭ[�r�          ��꺎^�g�>!ܙ	q����          dP�u�e�;��`���;w�\\�p!w          �F##�	`��T�|�r�>}:w          c`8�`0ȝ�{0pgjmnn�ɓ'sg          0F��~�F���w�R�׋n�u]�N         `�EUU����3u��at:w�          𮊢p��2pg��u�N'��ȝ         �K)EQ�Rʝ���35RJ���o��F�          &@]�Q�e��������+�ĕ+Wrg          0AF����1pg*�?>Ο?�;         �	4����� ܙ׮]�����3          �`�� �Ag��D��ڊ'N��          `
����F�3f��;�,�XYY���r�          0%ʲ�O�����4�bee%��a�          �HJ)ʲ���s��$w&N]ױ���^/w
          S���(�"RJ�Sf��;g}}=nܸ�;         �)f䞇�;����q�ҥ�          ̀������Θ)�L��/ƹs�rg          0C��a��3����p���8u�T�          fP�ߏ�p�;c&�3�n߾'N���R�          fTY�QUUg��X��������(w
          3�(���:w�T3pglUU�N'��~�          ��R�z�H)�N�Z�R���ƭ[�r�          �[RJQ���.1pg,mll����sg          �o��*ʲ̝1��;gϞ�.��          �w5���w��;c����q�̙�          ��a��S�������'O�̝          w����h4ʝ15��^/VWW����)          pO�����rgLw����tb8�N      ���w�Qr�w��ϯ�[]-ɹ !!�3��L�$1�L�,0���!��aM��K�f`�̲k�n�Ͱ1�d��rr�%`�d21��j�dɱ#Y�e˲eYr�/U��a%⛤�~��_�s�t�U�����\���   �(SSS{^ ���t���155U:          .Z�9���"�\:eY3p���s:t(�|���)          p�:����%2p��#G���ӧKg          ��i��133S:c�2p��'Nĉ'Jg          �����3r�H�,�ӧOǗ����          �hfggcvv�tƲc�Β�Ç��          �E733���3�w����t���F��.�          Kbzz::�N�e���%1??���177W:          �L�9&''�ܟ'w]�Ӊ����d�          Xr9瘚���s键g�΢�җ�gϞ-�          �t:#�����Eu���8u�T�          (��n���L錮f�΢9y�d?~�t          t�������-�ѵ�YgΜ�{ｷt          t�������/�ѕ�Ypq�С�9�N         ��455�v�tF�1pgA������W�          �s����N�S:����`嘟����ј��)�    �R�F�����#b��#��3]$�4�s������?��.���3\�'�����    �%�����k�FJ�tJW0pgA������~0    �2�R�<??�9���و����xjd>S9�1�R�N)=�s>�s�)���N�s���7�gfff&#"fffεZ�eqd�M7��������������^XUU�t:�)�zDDJ�)��s~Aι?"֦�.;�3k�q}D��گs���_cݒ��     �@�9&''c``��="�����}�ޟs�X��ݗ���8y�d�    �g3O�ϝ�����gs�g��:��t�UU�����v:��9�n��\�v"b�֭�#b}�V{aJ���N���s�/���"�E�?�0"^�5_��j    x.===Q�?ۛp��\�x ����    ��҉��9�ǫ�:}���rΏE�骪N��NG�����Gׯ_��k�/�Li�Vk�^��8����1������û�    K���/֬YS:�(w.ɩS����å3    ����"�dD�L)��9�L)=�s>�#�t__����N��r�ZV��n��E}}}���9�Dķ�_ZUշ䜿9"^O��    \�������-�Q��;��ٳ1::�N�t
    ���Ώ���S)��hD<��tN���#�����Z-O8�lm߾�%����/���F��RJ/�9�,"^v�{������    �2P�ף�gu����;err2���sss�S    �򞈧N]8"�朏VUu���<���s��/�6lhn��q�M7�h͚5��n�_�R�"�tE��[���Q+[	    ��R�z����{����6;;���1==]:    X|sq<"�Fă)���@��9��t���z��jy�P���[�v��SJ���oM)]�s~E��������p&    ��RJ100UU�NYR�\�N�###��O�N    �t�?}��ǡ���===Gϝ;w��j͗����n��E���W����t:W�����c�    xnUU���@��z������{w9x�`�>}�t    parJ����#�h��hUU_�|dpp�L�@`�|�#Y7==�_;|�9_�R�'�m�S�    ��Z-�����w�����{�w�}��C��     ��LD���SJ_=��^���k�/�t��~�����������"�����2����+��    Ϥ��'��z�%a������Ƒ#GJg     O9wG�WG�===G�����SJ�p�L�t�M/���"�tE��yMJ�ʈ�"����@�>    X����b͚5�3��;�����q��wG�~/    Kh>"�����N)L)z��'�k�Z����c�޽�cǎ}[�V{M��yMUU��9_������4    �"������[:cQ�����bdd$��v�    X�NF��)�C9�#�����p�՚,�LZ�V�^������_W��^WF�k��    M�^���������g455���177W:    V��)��N�`UUw������^{�x�0���j��֯_���)��Eĕ9��E���    `�X�vmTUU:cQ�����b���19�(    �H'#b_�y_D������M�6�,Pʞ={.���������_�s�*"��   ���R����9r7p��t:��뮻�ܹs�S    `9����"b�W>����S��[����˾����ʜ�k"�-���    ��UU�R�O�/H��kܗV�9>�>�h�    �FO�S#���H��������j͗X)r�i���WTU�Ɯ�"�)�7E�KJ�   @����z�^:cA���������    �=��UU���On�Z��] +ZJ)Gđ������n��-UU]W������Fċ�T   @w����������/��`���W�<y2���/��    ���xj̾/"�����]�՚.���ٽ{��N�ꈸ*"��9wD���    �y���5k֔�X�DDę3g����s.�    K�XD�MD|1"�X�ׇ�����I \�V�շnݺ�Gě����Q   �%P�ף���t�%3p'���bdd$��v�    X�qWJ�Έ�WU��7m�t�p Kd�֭�k���s�oK)]o����   �ŰF�����L���L�    X(�"�9�;#��Z�������Q t��{��N�8��U9�E��qe�.    X(k׮��Z�ojhྊ���ؿ��{�e    ���qgD|���;7m�t(��KG�|l۶�)�7WU����:�|UD���   ��QUU���e;r7p_�r�1::O<�D�    �s�ň�|D|~~~��o��s�� XaZ�V��u�ޔRz{����ֈX[�    ��Z��z=R�������b��q�=��#�<R:    ��|DܕR������n�?o��Rۻwo����o���#�mqMD��l    <�Z��3.���*t�ر8v�X�    x:s1z~�~G�V�sppp�t |��{��N�8�N���;#�Ņ�    �����F�b�ʜ:u*>\:    """�4�s��������������뮛)� ��jU�ׯ}���#�"��"��V   �S֬Y}}}�3�7�U�ܹsq�]wE��)�   ��Վ�����>11�V�5]:
 R�ժ֭[�Ɯ�5)�k"��X^�d   �����Gooo����}�����������+�   ��s4"�H)ݑR�������A ��v��U�t:W��v~���S8   �U$��z=j�Z��d�
������pLO;   �ŗs~,������V���M��N���u���UU}OUU�䜯���J7   ��b`` ��*���W�v�###166V:   ��k*">�R�����144t ��KG�r�}��o��kΟ�~MD��p    +TUU100)u{��3p�4�ӧO��    `�9w��������k��v�t ��V�Z�n�s��TU���["����   `Y���{wV}��w�}��C=T:   ��a:"��s�#��顡�C�� `5رc�7��ޑs�&"�/-�   ������z�t��2p_��?G�-�   ����S�����b˖-c�� `5ۻwo����op�;    ���/֬YS:����@�=�X:t(rΥS    X^�#�?��,���7o��t ��n��o�����������xQ�$    ��������-����0ccc122�v�t
    ����W)��{{{��뮻���A ��;��[RJ��9�7"^U�	   ��^�GOOO錯2p_A���cxx8fggK�    �ݎ��n�t:������ƍ�J k���W���w��~"�����J7   НRJ100U�O!��sss1<<SSS�S    �>��؟s�=��顡�}�� ���cǎoL)�H��]����t    ݥ�F��+@�Ӊ��+Ν;W:   ��1���O�j�Ooڴ�d�  ��]�v����۪�zw��'"�e��    �UU���@�Tvbn����СC��c��N   ��'"�OsΟ����O�Vk�t нZ�V500𖪪~,��c9��K7   PV�V�������ܑ#G��,�   @9g"�?�o������Vk�t �<�ڵ�5�v�'RJ?�U�   �2zzz�^�����2���ǽ��[:   ���xD�Y����.��/6n�8W: XY�2v��)�W��   `i�Y�&�������}�:s�L8p rΥS    X'�Q���j��K ��������zw��m�{    X�����ۻ��5p_����bdd$��v�    ��ɜ󧆆������ ���n��]�Z��"��#⍥{    X<)����������"��C3331<<333�S    Xg"�?�?>44��v �[�޽�����2����xU�    ���@�j�%����2�n�c���1>>^:   ��u."�4�|�e�]�7n�+ p!v����v��)�����(�   ��I)���@TU�4�[��\���ctt4�x��)    ,�鈸#�t����'[��d�  ���cǎ�RJ?�s�/-�   ����j100�$�2p_&��x�GJg    pi��ٔ�'����d˖-c��  �޽{kǏKD�/"~2"^P8	   �K����z}��c�;v,�;V:   ���sΟ��?��j�<S: `��Z��u���H��_���kJ7   p�z{{���Q�a���}��8t�P�    .PJ�xD�q����͛7)� �-v����N����"❱~g	   ��[�fM���-����ɢ�<p?{�l���F��)�   ��s."�4��񡡡Ϥ�r�  �n�u��着�SJ+J�    �����Goo�\���KMLL����c~~�t
    Ϯ�R�D���T�ٜ( �ܴZ�jݺuo���E�OG���I    <��R�����j���[����������)    <�C9���`��͏�� X)v��U�9�+�������%   ����b`` ��Z��.���j���������)    �#9�Ǫ���v���7o)� ���|�͗����LD�?"���9    �#UU���@��p�t�.s���8}�t�    �^'"�*���m���S��  V�;v\��*"��   �Z��z}�F��]��z�t    Oy8�􉪪nݴi���1  <��o~AOO�O��6朿�t    ===Q���Z�]���#G���    X���ٔҭccc�j��K ��v��qUJ�gs�?/.�   �����Ś5k.�:�]���C�Eιt
   �juo���z{{���?U: ��j��ׯ_���/G�;c�   `%Z�fM���]�5�����>p?w�\�u�]��tJ�    �6S�Ɉ��F��_RJN  Xv�������_�������t   �jS�ף����������ؿ��ΖN   XM��s�ݹ����Ї>�x�  G���[�~�{ϟ�~M�   ��"��z=j������,��:p������ᘚ�*�   �t"�r�{���nwZ; ��cǎW��~%�����t   �J�R��������vz�J�w:��'�|�t
   �Jw*���9��z�t  e�ٳ���ٟ��_��ו�   Xɪ�����H��&��>|8N�:U:   `%ۗRڳnݺ?޸q�\�  �ώ;���F�OEDo�   ��V���������;r�H<����3    V������G���h�  ��m۶�4��s)�_��o-�   �����F��~���z衇���+�   ��ܓR�3??�mٲe�t  �S���Y�~�{;��RJo/�   �����}u    IDATŚ5k��cܗș3g����s.�   �"����t:[���nO)y� ��m۶7TU�+񾈨��   X	�������9g����bdd$��v�   ��n&"�VU�upp���1  �l۷oID��)�D��K�    ,wQ�՞�1�lff&���cff�t
   �rv2�|���܇?��=^: �ե�j��_���9�FD|O�   ���F��n���pLLL�N   X������[��7n�8W:  v��quD\�}D��   XvRJ100UU=��/q�[���s����O<Q:   `�iGğw:��7o�|g�  x:۷o����6�9"^T�   `9��*֮]��g�H>�N�*�   ���Eĭ�v��-[��(  �Ǟ={.�������>"^Q�   `���j100�u�7p_ǎ�cǎ��    X.�9�v�V�388x�t  \��~������?�snF�kK�    ,��������g��N�:�.�   ���WUu����T�  X(;v�:"�DĻJ�    t�5k�D__�W�lྀΞ=�����tJ�    t���pD��+_��?ܰaC�t  ,��;w�1�)"�eD�J�    t��������311�������)    �(G�gr�{���K�  �Rڽ{��N��9��=    �&��z=j����B������ᘞ�.�   �mf#����j����ݥc  ��={�|���̵)�DċK�    t��R�_�v��������)    �d*��;���۷l�r�t  t��|�#�&''%�Ԉ�o.�   �-��2p�T���t   @�O)������-[�<\:  �ٞ={�����\D�ZD��t   @70p���w_<��C�3    ��XJ�ߥ���)  ��G?�������9������=    %�_��Ǐ�ѣGKg    �v:������[6m�t�t  ,g�V�Z�~��u:�SJ�.�   P���Ex���СC�s.�   Pʣ9�]n�Z��c  `%i�Z�ڵk�ED�۔қJ�    ,%�t�ܹ�뮻���N   (၈�]Uխ���S�c  `�۾}�5)�ߌ��)�   ��/���T���\�   ���@D������`�ƍ� �%�k׮�t:7F�?+�   ��ܟ����ؿLNz�m   `Uy4�kbb�Z��t�  X�Ο�~sD\U�   `1�?�N'FFF��'�,�   �drΏE��Z��gppp�t  ��r�iǎ�J)�o,�   ��zJt��s:tȸ   X-�9o����p���Vv  ЅRJ9">�s�}׮]?�s���xU�.   ��`���9�O�.�   ����?�n�w�p��J�   ������V�������X��7#�;Kw   \�T:��۷��9珕���?��{o�[   ,���G���yӦMgK�   ��jU��7E�w��   �������q�����-   ��H)MF�o��v�)�  ,�V�շ~��_�9�zD��t   ��0pccc122�v{)o   ��#������[�ly�t  �xZ���ڵk?�R�!"^X�   ��0p�G���cxx8fgg��    K���R��h�[:  X:�v�zq�ys�������   x6�_��n���pLLL,��    �DJ�Μ�CCC_(�  ��u��W�j�_��_��Z�   ��c�~^�9FGG�'�X�[   ,��SJ76��J�   �c��ݯn��7Fď�2��1   ��t��K5p?|�p�:uj�o   ��RJ�s����_��7l��.�  t��;w~o�ӹ9����-    _a���<���y   ��p:�c͚5�\w�u3�c  ��a���פ�vD��K�    ����#�<��s�b]   `)L�w�|�׎��  ���{��x���O)�FD��t   �z���ٳgctt4:��b\   `���d�yK�ټ�t  ��m߾}mD4SJ�#�^�   X}V��}rr2���c~~~�/   �����n޼���!  �ʳu��W�j�_��_���t   �z�ʁ���l����B^   `)<�R�����O��r�  `e۱cǛSJ;s��W�   XV�+���v����   ��D�������l47n  ����������GK�    +ߪ�:t(���Kg    <_���D���'�f��j��j  Xr�f����㯎��#�\�   `�J��˾}�ޟs��B\��{~x!.   ��RJ��t�f�`�  ����[�y~~�7"�"�V�   XYV������q��w�   ��)��h4>^:  ��l۶�UU}8"�.�   �U逥�裏����_:   �L����_e�  t�͛7�4��O)m��K�    +CO��v�ܹ��{"�\:   ��ܞs�nhhȫ� �e#��#��۷�YD4SJ7DĚ�Y   �2�J<�}���?�����٩��������   X(�E������t  ��ڹs�w�o��.�   ,OU��2770n   ��D��ƾ����  +E�Ѹwhh�Gr�c�{   ��gE����t⮻�s��-V   ����ɔR��h<X:  `��ڵ��n�����DD�   `yXq��s:t({���   �#�N�W7o�|g�  ���{��+����xO�   ��U��ѣG��  ���R��9߸~��f�  �6�6m::44�ޜ�{"��=   @w[Q��'Oƃzgo   ��ܞs���l�6n�8W:  ��f������+s�7F��?   �V*�\�������Ǟ�q�?�x8p`)�    ���SJ�s���x�  �n�s�����ψ���-   @wY'����šC�Jg    DḐ�����W�  <�F�qW��xkJ��"���=   @��)p����ctt4��v�   �����h|�t  @�K)����m�����m��M   @y�t�sٷo��s�{�������������Rg   |�s�\~���ǆ�
  �"�ܹ�9�ߎ��*�   �S��X�N'8`�   �v[�ݾrhh跌�  .^���lUUoL)�s�{   �2��	��S�N�H   ��x$����F�S�C   V�]�v�������xs�   `i-�܏=j�   �t����k��  ��������F���m�  `Yv'�?��#q�=��L   V�c��CCC��t  �j�m۶飯�w"��[   �ŷ�Np?{�l�{･3   ��'Gĭ�z�u��   Kk���G��;#bcD���   WO��krr2<�N�t
   ��|9��K�f�s�C   V��R��[�n�z{OOϿ�9��t   �8��	�3331::���S   ��c>��������   �a˖-7�M)m��ӥ{   ���J<�/|�������=>>^:   X=F��������+  �ӻ�[�y~~����[   ����'�?��W�   Kd.��o��ǯ2n  �n�_�����9矌��K�    ���N�   V�C�F��Z���1   <?�fsoOO�kRJ�o�   ��-��;   �b�q�����������  ��]����Ə��6D��{   ��g�   �f�r��|hhhc�՚,  ��i4�E�#⳥[   ��c�   �V����k6��+  ��z��h�3"6F�D�   ����    Xb����l~�t   �#��#��m۶}���ߏ��'   ϓ�  ��������  ��7o>2>>����1[�   xnNp   V�3)��h4n+  ��j�Z��u�Ν�s�DD��t   �̜�   �t�m�ۯ7n  X�������7���DD.�   <=w   `���9�x����[�l9Q:  ��Z��t���`�����x�t   ���  ������ۛ�fkÆ��1   t�͛7�e���9�?+�   �C�   �J�z��O��_�  �{5��G�����G�L�   �)=�    ȹ����l6��t   �CJ)G�om߾�3)�?��וn  ���	�   �J�_s�o4n  �b4�̓UU}OJiO�   X��  ��l>�|��_�}�f���1   ,_���S�F�9��!"/�   ���;   �\=�s���l�6l��.  ���l6���n�!��_J�   �jd�   ,G���껛��ߔ  `�ٲeˉW����9���=   ���   ��|������<S:  ��kÆ�f��J)�`D�*�   ���;   �\<�Rz{��l�Z-��  �$��g����"��[   `50p   ��۫�zC�����!   �>[�l91>>�����E�   ���  �n6�s�q||�����gJ�   �z�Z��f���9�wq�t   �T�   @�:��t~��l�Z����   �
�f�v����ҝ�[   `%2p   ��===oڼy��    ]g˖-'���~ �|cDxQ6   ,���    _����hܔRʥc   ���Z���h�ܹs8���xA�&   X	��   t�3�/����w�v   ��F��UU�)"�n  ����   �#�Z��CCC��t   \����/����D���-   ���   E���h||�m�6m:Z�   .ֵ�^;>44���1"�J�   �re�   �2�s���h��V�5Y:   ���ЭqMD�*�   ˑ�;   ��rΏ��~��ln-�   mhh���v�M�7�[   `�1p   �TJ��N��F����-   �X�l�r������[   `91p   �ҭccc�|˖-�  ��v�u���RJ��"b�t   ,�   �R��9������V�5[:   �R���x����H�   �v�   �b{<��C�f�c�C   ��f��_��zS���J�   @73p   ӁZ���f����!   P����CߗR���-   Э�  �E�s������7m�t�t   t�V�5=88�39�"�S�   ���;   ��RJ{&&&�}�u�=Y�   �MJ)7�ͭ)��J)M��  �nb�   ,�����5��Z-��  ��h4�������n  �na�   ,��UU}���x�   X.6o�<RU��F�ߔn  �n`�   ,���������!   ��lڴ�d__��s�^4  ��g�   \�OVU��n��۩  �E���f���ޟR���ȥ{   �w����{�����;�}�9s撹$3�ҖD[��ZZW��]�
4���ea�A��beDN����s&Ѷ?�1%�(�Z,ڸl23ɀ EK-�*��B��䜁䜽O��A��df�콟}y��J���{���}>�9  ����^�����n����-   0�RJ��������@�   (��   ؊AJ�Ǫ���i��t   ̒��5��Ԉ���-   0n�   ��:�s����^_:   fU�����N�["�K�   �8�   �/"�^�wG�   �u�n�O666�%��[�[   `\�  �����-u]���!   0/n��ϯ��=-"�U�   ���   8w/,,<���O�  �y�4�UU='����-   0j�   ���yϞ=O?|���+   �*��{�^/��A�   w   �lrD����^p�С��1   @D]ׯ��g���X�   F��   8�AJ�Eu]ߘRʥc   ��Q��{ڶ}jD|�t   ��;   �p���SU�K�    g���~;"�ED|�t   ��;   ���#⻪����!   �����"�I���-   0,�   �i�m�������   �O]ן�t:�*�   �`�   DD|"��/VVV~�t   pa���9�E�]�[   �b�   ���t�TU��   ����Z__��xW�   ��   0�>���qU���t�   ��4M�QU�s"�ե[   `��  `~���t�z�7|�t   0)�\�u7�|�t   l��;   ̡��[��ׯ�v�_*�   _�׻%����ȥ[   �B�  ����S�N�p�4��!   ���z����k"�w    L���   �X���������   s���w��U�����J�   ����   �DJ閺�̸   �KUU�J)]�n  �s1p  �9�Rj��:R�   (���_�t:�_*�   ���   f[��nUU/+   ���vo����-   p6�   0�r�y���W�   &C]׿�*"�-�   gb�   �i�RzA�����!   �d�����m�m�W�[   ���  `�lD��WU���!   �dZYY��N��Ԉ�l�   �j�   0[6#��u]�j�   `�u���5����(�   ��  ��䜟_��{J�    �auu����_F�gJ�   @��;   ̊AD\���n+   L���ՏG��;   ��   �� "~���_.   L����0���#�J�   0��  `�RJ?T��;J�    ӭ��}4�����|�   旁;   L�6"~�����   fCUU��m[#w   �1p  ���F��~[�   `����|�G���n  `��  ���)��u���!   �lZYY�HJ��  ��3p  ��#�UU��t   0۪���N����-   �w   �.����t   0����䜟�J�   0�  `z�ۺ�_U:   �/�^�期�n  `��  �H)���룥;   �����ND��GD�t   ���   &ߛ���KKG    �����~$"��-   �.w   �l���+�MJ)�   ���9��Jw   0��  `B���---�����[    N��z?�RjJw   0��  `��~�m۫���,�   �pUU�,"~�t   ���   &�������z�S�C    Φ��ՔқJw   0[�  `������3VWW�J�    <��R��+^�R�  ��a�   ����~�;n��ϗ   8�ٳ�q�t   ���   &�r��8r���-   p!:��������H�   ���;   ���R��^����!    [���|�`0����d�   ���;   �զ��WU�ݥC    .����G�3"���-   L/w   (�[Uկ��    ���� �����K�   0��  ����-u]��t   �0�z��n���#bP�  ��c�   eܶ��vC�   �Q��zw���-�  ��1p  ��;����CMӴ�C    F���7F��Kw   0]�  `�>��������K�    �ZUU7D��Jw   0=�  `|�"��������   ��R޳gϏD�=�[   ��   0_�t:Ϭ���J�    �ӡC�6;���E��n  `��  ����w���)   PB�۽w0|WD�W�  ��f�   #�s����w��    (iuu���̈�(�  ��2p  ��zK�׻�t   �$���7SJ/*�  ��2p  ������ҡ�    ����_�9�Z�  ��d�   ��KKKW///?X:   `Ҝ:u��R�O�;   �<�   0|�w:��Z^^�\�   �I�4M�cǎ�E��,�  �d1p  ����9o�����!    ���k�]ψ�O�n  `r�  �p����(   0VWW�<����x�t   ���   ��mu]�l�   �iRUՇRJ/,�  �d0p  ����N�P�   �iTU�[#��;   (��   .�g��ww��/�   �V{��YN)��t   e�  ���w:�g���~�t   �4;t���`08�.�  @9�   pq��n�}�#    f����gRJϊ�K�   P��;   lV��    IDATQ���u]�t�   �YRUՇRJו�   �w   ؚ��:u�P�   �YTU�SJo*�  ���  ���|���i�X:   `V�޽�ڔ��Kw   0^�   pa)����zZ:   `�:th3�����l�   ���   .̿���d�   �y��v?�s����n  `<�  ���}�W�R:   `��z����n*�  �x�  �������s<�0   �1[[[�)�t�t   �g�   ��o�����?W:   `5MӶm{MD�y�   F��   �!�|�����Kw    ̳^����N�"�_�  �a�   �(rοQ��+Kw    ��v�M�   F��   ���RJ?�RʥC    ������#��   ���;   ��f۶ϩ���J�    �7��i������O�n  `��  ��VWVV~�t    �������ҳ"b�t   �e�   ���UU��t    gWUՇ"���   ��;   |����ڶ�єR.�   ��[__�9"�[�  ��1p  ���;��VVV>S:   �sk��M)=?"�+�  �p�  �_K)����_/�   ������"�%�;   w   ��?H)���    ���u����;Kw   p��   ���m���v�T:   �����|qD|�t   ��   "~|ee�#�#    غ#G�|�m��EĠt   [g�  �\�9�o}}�ե;    �x+++��s~y�   ���  �yv�`0x~�4m�    ��ԩSMD|�t   [c�  ��J)��#G�o�    ��i�~�ӹ&"�K�   p��  �K9�WU�k�;    �n��'�Z�  �g�  �<�����u�#    ���~.�t�t   ��  �ytm�۽�t    ��RʝN�PD��n  ���  0Wr�o���ݥ;    �Ç""���   ���  0O>���p]�    Ƨ������;   8?�   ̓k��#    ��R^XXxaD��n  ���  �9��u���    ���Ç?�R��t   �f�  �<�����u�#    (����lD/�  ��3p  `\��v�-   @9)�����X+�  ���  0�RJ���ݥ;    (���ßH)]_�  ��3p  `��۶���    L���������   ���  �Y9�^����;    �MӴ9�C�Y�  �G2p  `V}���_*   ����z��R��t   �d�  �,ڈ�C)�\:   �ɔRzYD���   <��;   ��u]�A�    &W���R�ӹ�t   e�  ����N�ss�    &_�۽3"n/�  ��0p  `ּ���~�t    ӡm��"����   ���  �%���x�    �����g"��Kw   �e�   ̊/,,,�JG    0}����,�  ��;   �c����Q:   ���4M�s~QD�K�   �;w   �^J�w����t    ӫ��}4����;   杁;   �.��6MӖ   `�mll49�ϕ�   �g�   L����VVV�_�   ��w������t�m�  �yf�  �4[o����    ̎���7�?\�  `^�  0�r�GWWW��t    ��i����\�t  �<2p  `Z���۷��t    ����FĻJw   �#w   �RJ������    `6�^D�*�  0o�  �Fǫ����    ̮���O��n)�  0o�  �6���%�#    �}kkk?Z�  `��  0m~zuu��#    �}M�<u�  �yb�  �4�����\:   ��Q���#��;   慁;   S#�t����[�   ���s�#"��   ��   L�On۶���#    �?�^�SJ�)�  0�  �
)��X^^~�t    s�HDl��   �u�   L�������t    󫪪?�9�R�  �Yg�  �4Xi��-   ���w�V:  `��  0��[��]�#    ����eD��t  �,3p  `�刨KG    �i;w�%">[�  `V�  0�n������    �Ӯ��������   ���  �I������#    ��������t  �,2p  `"�������t    <\�4��   ���  �I��R��t    �͕W^�Έ���   ���  �I����?Y:    �������8Z�  `��  0i//    �r�Wޖs�X�  �Yb�  �DI)�iuu�S�;    �\��  0|�   L����-�#    �|�:u궈���   ���  ���R�y��   0M��is�?Y�  `V�  0)H)��t    \�S�N���t  �,0p  `"�����v?]�    .T�4mJ�-�   C`�  �$x ����    �Ukkk�-�  0��  (.���no   `���-�7��   �v�   ���s��t    \�+���W#�OJw   L3w   J����O��    ��u���AJ�e   ��  ��ڶ�?    f������ϔ�   �V�   �s��������    �ai�恈x}�  �ie�  @1�(�     ö�����X+�  0��  (�u�����    �a����_(�  0��  (��    `T����Q�  `��  P������t    �����rη��   �6�   �]���MӴ�;    `�_�  � �   �U��s�N�z[�    �Ç,"�K�  �ib�  �X��o���    0�^z�{J7   Lw   �jcc����Q�    ��	_���l�_�  �/w   Ʀ��G۶����n   �Q�뮻�#�y�嗗N  ��   �������\����J�    ��m[XxiD�<�,,�:  �|�  0m�F۶����>���=�d    ��>��=)�E�N'\vY�$  ��`�  �X|����s^-�    #�����"�������<�`  ��0p  `�r��������i���   �����?�-r^��۱}{�ݳ�T  ��0p  `��0n?me�    0�_���"⊇��c��  pN�   ������~��o����    ��sN9��L?۷wol߾}�I   S��  �����Ѷ�Y޶��    �����p��?���1�   Lw   F�Qno?��G���q�    ��uRZy��ؿ?:s  ���	  ��i�6���^�������   �Qz�O���h�Y\\�K��W  ��1p  `d������G����l   �Q�7���.?p`�)   S��  �����<ߗ�����Q�    �(�<~��Gķ��k���۷oq  �t2p  `$��~�/�-���   ��J����ؿD!   ���  ��������~e-    0J�=q�["�__�{\vوj   ���;   #���{D���y��[    `�r��.�=KKK�wϞQ�   L5w   �nsss�o��CL   �����ۿm+����!�   L?w   ��"�?�w    �E��q��t߾X\Xf  ��3p  `�ڶ��m/��#�Ȑr    `d���o���m��)�8���   ���;   Cu������G���a<    Fe!�.��80�  ��a�  �P���a<f����A    0
�;���ԋ}Ύ;b׮]�H  �	�   �`0����#M���a=    �)u:G�����^:�G  L=w   �fsss��[����   `��gD�S����.�lX�  �z�   M���#��4�?�C   `���餶��K۶Şݻ��H  ��e�  �P����RD�r   �����O~~D|Ӱ��w  �/3p  `(���}U�4�>��   ��:y�䎔��F����틔�(  0U�  �h9�����<�M��   @Qy0X�W��ً���wϞQ<  `�   p�F<n���Ɣ�sG}    �������:��<�K/��  ���;   m��9�|뭷��A    p�����g\�o_t:�  �|�  ���s��`0�������q    _�������v��,,,ľ�{G}  �D3p  �lnn���7M3�[�    ��R��;�q���.�1   ��  ������y�eq�8   `��s�=�8Rz��ۻgOt:�  ���  �-�9G۶�>v���n���>   �����5i���N�{���q   ��  �-���m?]�`    ��=Ǐ������}{���H  ��a�  ���RG[�4�Y�p    f�?���)�[J�}�}�R*q4  @q�   lY��O{��^���%    �]_�⑈��g/..��K.)q4  @q�   lI�q{D���w�}/-   ��y�]w]uɆ}{��<  �w   �d0�N���O4M�wJw    0[څ�[sĮ����W�x  �b�  ؒ	��="bwD���    ̎�Ǐ?)"��t����c��3   ���  �6"�\:�k��yR�    ���߾)�LD��-nq  擁;   lBno?-E�k���   ��r����"���8��K/-�   0v~�  ���D�JG    0�����)���_m�Ν�m۶�   ce�  �i�6ڶ-�q&�4M���    L�틋����;n�=�   ���  �2�����?"^Y:   ����'��� �yc�  ����{D�5M�<�t    ����o_��7DD*�r&�  ��1p  ��L��="�皦�Q:   ��p���Gr�ח�8����صkW�  ��1p  ���9��8�'D��#    �|�;v����Kw��>��  s��  ��6�����4��޺   �dh;������k�{� �9b�  �y����RD�!"R�    &�=Ǐ??"�V��|���tL<  ����   �m��On��KG    0y������~�t��J)ŞݻKg   ���;   ���N؊�j�汥#    �,K��S����={J'   ���;   �e�no?mD��t    �����OI)�P��w���	   ca�  �y���#"~�i��KG    P�wܱ+"��t˅ڱ}{,m�V:  `��  8��s�Kg\�7�|�͏)   @Y�����H�	�;�j��ݥ   F��  �s�.�c666^]:   �r�9v쉑�;.��;  0�  8��GD<�i��KG    0~w�qǮ�қӔ�$v_rI�  ����n   �ǌ�#"^�4���    ��%�v�<RzB鎋�sǎXXX(�  0R�   �S۶���q��    ��=ǎ=1r��tǰ��  �u�   <������6Msu�    F�;�ؕRzs��}��;  0�f�   ����K'��뛦�_:   �Ѻd׮�GJO(�1L�  ��3p  �Q������ז�    `t�9v쉑�;��K.�N��  �]>�   �ڶ-�0*�k����    �ɓ'w�N�-iw)�صkW�  ����r   ό����~��ѣW��    `���D�ו��ݗ\R:  `d�  8�9�_�����4���    3�w��=�#�;F��  �e~�  �Y���="⪈xi�    .ޱc��N��M�;F�]�J'   ���;   gնm�q��i�o*   ��5M����%"�n����XZZ*�  0�   �Q�9rΥ3�e{D���[o�Y:   �����O�F��Jw��[� �Ye�  ���	������-�#    �p'��E�7���];��   �&w   Ψm��	%�X�4�Y:   ��w������Έ�Q�e�v��  �Q�   �����"���y\�    ��`�ʈ�����w  `V�  pFsz�{D�c#�M��;    ���/.�Q���b,--��   :w   !�9��%}g�4ו�    ��~��;�v�xK��E���U:  `��  x��`P:a��i�o-   �#5M�l������7�v��Y:  `��  x��mK'L�mq��7�|�t    u��xc���Jw����  �2p  �ܿ⊍����3�    ����~j�t�t�$p�;  0��  x��`P:a�|G�4U�    "N�<��N���-�`qq1Kg   ��;   ��s.�0i�C�4O*   0�N�<������-�d��   ���  ��h۶t�$Z��_n����!    s�mo��'�Θ4;�o/�   0T�   <���Y=>"��4���    c�޻�~z�y�t�$ڱsg�  ���Ky   ���Q=="�"   `�N�<����[����ܱ�t  �P��  �C���M7�x�U�#    ���?��m�����n�T;� �c�  �C���b۶�v�M7���!    ���/|�U��KwL�m�����P:  `h�  x��r`0�Z�4�J�    ̪�'N</�����`�[� �b�  �W�_�o��7��    �E�;~����^Λ�;  0K�  �
����i~�t   �,9q�ā6�_��z�y�n�  �w   ���}K^}�7^U:   `�<yrq!�W#��n�&np  f��;   _�s.�0�۶}W�4�/   0��`�xJ�i�}i�t  ���  �np߲����[o�Y:   `Z�<q�y9b�t�4Z2p  f��;   _a�~Q�����c�   �it�رoJ�[٢�R,m�V:  `(�  ���s�iwM�4/.   0MN�8q :�w�]�[����� �?{wg�Y�y�w�s�zɂi�HԠ����0"�+��ڑ	*�;h!I_�hDsCD0�0����0@c��ZN�4-jp'6LF��Nz���ι�
!饪���߯W?�<�Wu����� �"�  �������SkG    �����fJ��n�w.�  ���  ����v���HD�{۶m��   ���ݴ����'���\p  ��;   a����v�;_��W�S;   �W������+jw
� �Aa�  @DD�Rj'��-..���np:   ��LN>-Jye�A�;  0(�  ��W�>x��Ԏ    �%7ON>6��gѬ�2H֍��N   X�   D���*�Ŝ�o֎    ����)�/"N��2hFFF"�T;  ���  ���	���cccϨ   PӾ}�6t[��F���[QJ)FGFjg   �2w   "��}�5J);r��_;   ��RJZ��{k����*1p  ��;   ��kcCD�7��-�C    ������E�3kw:w  `�  `�v΋����5�9�v   �ZiOM=�D��v�0i�j'   �2w   ����N&�=v���n��u�C    V�����Sěkw� �A`�   k�I|[D��!    �eff�q�R�W"Fk����  � 0p  ��:.�9��v   �j�yb�a���@D�^�e���  w   ��R;aX�tll�ŵ#    VR��>��l~0"R�eظ�  w   �+*�\�s���    +a߾}R�����-�h��   �   ��Ո�cccO�   p*��Ǜss�,���2�FFFj'   �2w   ��-��;��]�C    N�9�6�>"~�v�0K)E�٬�  pJ�  �n�[;��EĮ뮻���!    '�=9�#�E�;�i�j'   �w  5Xj.    IDAT �߼���9�M�C    �W{z�y����|Qkd�v  �)1p  r���	|��|�k^sF�   ��gz�Qʛjw�e�f�v  �)1p  r�=���;������!    _O{jꩥ�?��V����0  ���   �MO���o��;�  ���gj�#���v_��  �w�j   �w]|�����=�   =cff�K�_D�i�[�Z͖��  @�9  ��+��N��=+"��v   �ͻw?"u�qV���  @��T  0����/圯�   ��'&��6��[���f�  �Sb�   ��Ws�/�   ����s���dD|k���  @��T  0�\p�+����   �p���|�h�ySD|G�X��  �s�j   ���{)������sjw    �a�޽g�"&"Ⱶ[8>�V�v  �)1p  r�}�QJyk����!   �`۹s�ƥ���GJ?P����;  ��<�   9��Ԉ�����]V;   L;w��x������i6��   N��;   ��f)�m9�g�   ˿�?�v'�w  ��y�  ��Ռ��666���!   �`عs��36l���}+�T;  ���  @k�R�>66vi�   ���۷o��7��D<�v'ϼ  �w�   �����?�9?�v   Пv�ڵnan�]Q�Sj�pj\p  ���;  ��+��N`e4#�9矮   ����������n���  ���   �HD��   �k|||��M�����;  ���  `��Dğ��v   ������s�:�G�E�[X9�  @�3p  ��3�cccϩ   ���;wn�N��%����   ���;  ��+��N`u4K)o{Q�   ������O߰��#�[X��9  п<�   ��J����9�j�   �7���o�Ng2"�T�   ;   ��_����!   @]�F��'"���-�.� �~�   ��X�y{�   ��v����Vk:"��v   �w   [r�o�/^u   �����Ccy��(�1�[X���	   '��   �ˋr�o�9�L    ���k��'Rzx�   8��  r)9�=�^4>>ެ   �����wv��["�a�[X[.�  ���  `���kh������s���o�   �������և"�k�����n�  ��f�   ��>���۷?�v   �r�LM=)5�Q�9�[   �D�  ��R��z�����뮻�57    {���Q"v��3k�P�76  ���   x����-�x�+Q;   8y3SS/�����v��  ���   ��xX�ӹe۶m��   ���������`��  �΃-   �o����~hll�Gj�    �g||�ٞ�|S���v���  �w�   C.�T;��rz)eg���j�    �o|||��M�vDJ�R���Q���	   ���   �j�"���9_Q;   �o�v��s�:kgD�|�zK)n�  ���   �/͈����յC   ��411qnt:{JJ?Z����u�  �s�   C.�T;�ޕ"�9��x�#�c   ��v����fsoD<�v��c�  �9w  �!g��q��|p����   �l���F����-��N�S;  ���   ��)���{s��   è=5�s%b&"ή�Bo��  �9w  �!�;'�1�m۶y:   ����ԋKğE���-�>� �~g�  0��9A�u��=9�j�   ��o�LO�1"^�|��q2p  ��`   �D���9��v   �v�}�9�6�/��_j��_:�n�  �Sb�  0�\p�$5#��sί�9�|   VЇn�����O��B�q�  �w��  r+#�9���C   `�'&�m�>R"��v���;  ���  ���;+��#b�u�]w~�   �g333?�������n���  �;w   `%<vyy�#۶m���!   Џ�SS/N���Kę�[�o�  @�3p  r.�������~(����!   �/v�ڵnfr��h���u���	   ���   XI�#�9��9g�;   ��h��goX�n"��K�[��˵   N�/�  �F��!+*EĖ��k_{Z�   �ESSS����D)O���`YZZ��   pJ,   ��򳳳�����o�   �dfr�i��["��j�0XJ)��tjg   �w   \pg5}����9��   ��RR{zzK���qf����  � �`    RJ�lgG����C   ��v��~���;����w�������	   ��C3   u����9���1   ��&''��ވxv�ۢ�  � 0p  ����tED̼�<�v   ���ݻ��J�#�q�[|K.�  ��   w�څKKK��_;   V�����ј��o���pX6p  ��;   �hx<d�}SD�<66��v   ��v�}z{jj<E�#�{�  � �`    ji�R���$缱v   ���w�~Dt��k�0|���j'   �2w   \p��gEć_�W<�v   ����ɧu���RS����;  0,   �^�:�����v   ��RJjOOo����P��ᵰ�X;  ���  ������ƶDD�   �c׮]g~O��=��ʖ��j'   �2�   D��;=�YJٞs~_�yS�   �?���߳at�o#�k����b�Rjg   �2�   """%��)G���9?�v   ܗ���˛���^�""]o  D�v    ��wz��qs����-�ܭ   {��=c�رSJ���M/YXX��   �"�   ���Y�����9o�  �p���z����GRJ��n�����X;  `E�  .���.����m۶�  �p������7%�Q�[�,�  �z  ��0p�/<���~hlllKDx�    k��n��gzzGJ��%bc��z\p  ��   _���0=�UJٞs~�_��j�   0�n��� :���R~�v<� �Aa�  ����N������n۶��j�   0�f&'//)������b�  �   ��w��ú�so֎  `0LNN>hfr�)������{�x�  ���  �/1p��"b����'s��R;  ��6==����>�R��v��w  `��  �%ͦ#���'E�m9�g�  �����7���[�썈o��'j~~�v  ��1p  �K����Eğ����׾���1   ���ɇ��i�L��="Fj���8f�  �   ����q����9��  @o����ّ��G����-p*j'   ��V�    zK�шn�[;N�wF�Grί��m9g�  ��}��mX���^"�,�c`��  ��   �
)��	�RF"bkD��9S�   zC{���]���X���v�����X^^��  �b�  �
��GE�S"����=�v   �����-�h싈G��z;  0hZ�   �-�f3���jg�J;���ޜ�"�Wr�k  �v����E��(�k��J�7p  ��|   |�p�#ⶱ����  `m�LN^���E��n����;  0h\p  �+��j'�j;���3�����9磵�   Xy�v�!��9".����w  `�8�  �WH)�3RD\�s���1   ��=�ӛ�ӹ-��.�  ��w   �F�шN�S;���"��s~æM�~��+�\�  �ɻ�[�Z^X��Rʳj��ZX^^�����   +�w   �F�٬� k�W<x�9��  ���3=�����"¸��177W;  `Ź�  ��h4�>4C���9籈�휳�g   }`׮]gn}m)��-�����   ��,   ���шxeD��;  @��������D�3�f]p  ��   |��R����R;j�������nڴi�W^�P;  �/k��ߐ:�ה�痈T�jq�  DN�  �5RJ���l9x��G�m���c   �����E�����Wۍ�Z��˱��X;  `Ź�  �}j4��tjg@/xt��ݗs~KD�z��h�   �a411q�H��;qY����  ��9>   �S�٬� ��_��w9�֎  6{��7�6��R2n�577W;  `U��  �}j4�N4܇�E���Dį��  d���:��K)?]�zͬ�;  0��   �O)�H)�΀^�"Ⲉ�mll��c   Q)%�LM]�m�>��p���   �*�  �O)%W����WJyO��Os��  0(����gf��"n,g��^�������3   V��   _��;�gF�'���^<>>ެ  Яn��֑����f�Ǣ�'��^�z;  0�,   ���M[]8N*��n����m۶�  �o����Ƚ�~,J��k�@�;:;[;  `մj   л��}O��ݗs~��޲eˑ�A   �즛nڴ��zu)���j�@�8z�h�  �U�;   _WJ)��p�Zq�c�>�s���1   ����f&'/_�j��qE��q+����\�  �Uc�   ��r�N�7EĻr�;���o�  �+���y���TJ��qv��7sǎE�ۭ�  �j�  �_.��)�hyyy�9�x�#�c   jٷo߆��dnF�]�xr��WG���   ���   �_.�Ê�[8�W9��׎  Xk{��bqn�HikD�������l�  �Uժ   @ok4�R�RJ�����9�?o�Z�~��W�v  �jj���R��_UJ��v�Y� ��;   �wXQ)"6///<�o��� ���o߾������)%�vX!�������   XU�   < wX�E�փ�]���k�   ��=��/���}��5"6��Artv�v  ��k�   ���êzdD|0�����sΟ��  pRn޽�%�וR~�v�#G��N   Xu�   <�F��`\O�9�vDl�9��  8��6/��҈XW���  �0�P   ิZ~G�������/�  �@�LO_����)m�vXU����X;  `�Y'   p\��f,//�΀aq~D�=�|i����k����k  �{�ݻ�Sj4^_J���-0,�9R;  `M�  p\��f�F?��v4�cdd�%/���  �v�}v�t�)/*>,�5t��  �   �F�)�(��N�aӈ�˖����s�݈؞s��  �}��mX8v���鼬D�Y��M)%�=Z;  `M4j   �?Z-�'�[#������*�   C����LOo^����l7n�:���F�ө�  �&�  8n��Ώ���?�m۶k�   �kzz���LM�RJ��o����ȑ#�   ֌e   ǭ�l�N ������-9�?o6�[���;j  ��扉�;��+S)ώ��=
z��Gk'   �w   NH�шn�[;���;��E9��#b{��7�  �Ii�ۧ���otSڒ"����hyy9fggkg   ��F�    �K��w��m���G�ccc[n��u��  ��q뭷����^��?FJ[øz��� �!c�  �	1p��vv)e���o�9_1>>ެ  ��RJ�3=���=�쏈7D)��n�֑#Gj'   �)w   NH�ш�R���=4"nܿ�����6׎  zO{j�{�����2)=�v��2p  ���{   ��V�KKK�3���R�x����Ҝ���A  @]�ݻ�7���Q�Sj� �رc���X;  `M�  pͦ�;��#▜�"��sη�  ������6KyY7�y�o��>q�C�   ֜�;   '��l�N N�E��9�F�X��s��  ���n�ώN�7��_-�R� ���  ���  ��R�f��N�v
p�ZqED<+���u����o��o�S;
  XY�v�:súu/�N��"��=��[\\��c�jg   �9w   N��Ȉ�;���"�eW�?"���  ������F���E�oE)�X�8y��  êQ;   ���l6k' +�����9��۷?�v  p����Gg���m6�OD�."�ۡ��  ��w   NJJ)�Ft���)���[����k��6l��-[��  ܿ���ѳ7m��F���M�{����t���l�  �*\p  ऍ���N Vރ#b�c�>966�����P;  �Z��z�������n���q�q;�C�G)�v  @�   ��Vˋ�`��SJ�~���O���m�9��  D�{��7���)�����P�	Xy��{o�  �j�  8i)�h4<Z;���=">166��o�ѫ  ��������R�x����M���v�q�ȑ�   դ�dǎo9p��skw   p�cqq�v�v>�R���3�x�UW]u�v  �����9�6=3"^��V߽��'︣v  @5�   ��n�sss�3�����xSD\�s>\;  ͭ��:r��{.M)�,"��v�v�������S;  �w   N���\t���@wE��G��r��֎ �~7>>>z�Yg=3E\)=�v����n|��|�  �V�    �_�Պ����@gG�ֈ�*��ƈ�����M  �wv�ڵn���sR�5�-�{�:�=tȸ  z�   ����w����/�9�uddd��_����  �׵��ӣ�yn|��������^/G  0p  ������lF�ө��wzD\�������[���\}���\;
  z�޽{�XZXxa�t~�Dl��Է�����  P��;   +���*#�W���_�s��F��k����kG @m�v�!��xy~��qf��{�R�T   0p  `E������b����F�e�n��9翈��眧jG �Z�����f)W�N������jｷv  @O0p  `E��\q�O���"⢜�G#�G=�Q;.��?4  h333��N�ũ�_(��=@oZZZ�#G���   �	�v�ٱc�[8���   <����XXX���O��~�3�x�UW]u�v  ��RJ�yf�Rʕ���=@��_��~�s�3   z��;   +��ѣ����xSDܐs>X;  N������g��̔�oFģk� ����sss�3   zB�v    ���lF�ө���s#bkD\�s~s��z��W_���Q  p����{����/G�oDķ�����q;  ���;   +jyy9���kg ���"��9��1  �����o�N翦�痈3k� ��sā;יִ  �3\p  `E�Z�H)E)�v
пqQD\�s�hD�p�y���^����]  333��N����\-O���*��]��   �).�  ��bi�XQ���#�9�j�  0|���G�}���^J������=�`��С��w��   �)�   ��n�sss�3������9��j�  0�>�k�9�u�~9JyQD�_�,��㎸�С�   =�U;   ���h4��hD�ۭ��uqYD\�s�pJ��\p�{.��N�0  ����#[/�F</J�X�<���q����   =��  �U1::���3��va)������ﱱ��+��q��2  ���sn<�	OxrD�8"�V����@�����(���   �9�   ��V�)%_�k�;J)o��W����h���k��X�(  ��M7ݴi]��KQʯD��k� �ᮻﮝ   Г�  X5�V+���jg �㌈����^�s�hD���3��㫮��X�0  z����������1�����8:;��3   zR�B�cǎ�8p๵;   8q�n7���jg ������a��+    IDAT�*�  �v�ڵn�u?U��GJ���ӧ>������   =�w   VM�шF��n�v
0�΍�-��LJ��\p�{.��N�0  �V��~xt:ϋ��R�Z;PK�ۍ{v  @���Om\p  �oKKK��u�@o�dJ�K)�s��v  �'��x����xqD<-���Q`���]wŧ?���   =��?�1p  ����QJ�����#��)�?ںu랈��
 `@LOOs��_.Ϗ��k� �{�?�86?_;  �g�j   0�Z�V,--�� �j�#�Y��g�?7�?]� ��0>>�<gӦ'E�Q�3��B�t���v  ���;   �������3 �G7"fRJo.�����r�   ����w[�_H���D<�v����;�C���   �i�   ��RJ�l6����Nx ��xj)�q ���f����\s�'k� �e�v�Z�qݺ�*�\эxJ��J�(����h�  p\p  `M,//Ǽ�/��?�9�U� Z7ON^�M�9�܈8�v�����}.>��/��   �y.�  �&Z�V���7���ӈ���ϫr�;��;���ڏV� 
{��=cia���}^7���p2��n�u�`�  ����;   kfii)jg ���G�xD����*�  ��s�^����e%�"���M �⮻���gjg   �w   ��ѣGk' ��nD�eD�#"ޙs�� �$�'&�3�gFJω�o���R>~��177W;  �/�j   0\FFFbii�v�JjDą���9��E�;r��Q�� �[n�嬥��ͩ��#�k� ��#G��  � w   ֔�;0�Ό��"Ⲝ�g#bG����k����T� �)����>��?VJ������1��_>pR�宻j'   �����hǎo9p��skw   �r�;�N�v�Z)�/"�9::�����e�R; �����H��e�̈xp��ն���k���   }��  �5��t�رc�3 j�D�G"��ׯ�������j ���''/�F�|J�����= k�ӟ���   '�U;   ���l6��hD�ۭ��֚qaD\8??C�y2"�u�i���%/y�l�6 �s�����f�g���ݔ.���km ����r�}�`�  ���;   U,//���|��^q,">�R��R�D�y�v ���馛6�6���.���D|	���������w��   �;.�  PE�Պ�R��@Dl��ͥ��qO��)�w]p��.��N�8 ��grr�A͈���6GďE�H�&�^��t⮻ﮝ  Зz�j��   �kii)jg ���F�{�Ɵw��眻��  v�ܹ���,��dD����k���ⳟ�\�  ��d�  @U�������"�)�w=�!��/x�R�  `x���)�nwsJ�#��M ����}�㱸�X;  �/�  P���/� N������һJ)9g?H��n��!u�?��v/N)�LD�V�	��u���O��L�  ��ժ   �p5p8q�"�R�eqo�ygJi�ƍw��%/�� ��[n�嬥���SJ�S��%b4�����S�����   ��z��(�  ���B,--�� �㋗�߽q�ƛ����155��F)OK)m������M ��СC�w�Q;  ����  @u���� +�̈���r����|�yoJ��f�ϯ���� ����oov�?U��G)O����� ��v  @�s�  ����;����j4;���ڿ��R; X[333�N���H颈x\��As��������   }��  ��PJ����� ��S�;��R�D�y�v �������t��"..?�\�	`�}���cnn�v  @�3p  �g��P�=1X�~��^�җ� ������Rzr�۽����Kę�� �����'︣v  �@h�   �3::j���Ί���y~~~1�|KJ郥���׎ �͓����JJG��K)͔R��a C��w�Y;  ``��  @Oq���|>"&SJ;׭[��uw �;w��x���O���Gķ�nf��p�  `Ÿ�  @Oq���<$".+�\6??��s����Δ�Ե�^����Z����������#�G"b��z���  V��;   =%�������X;��Ԋ�K)�R"�|gD�v� V�+� ���C�bvn�v  �@1p  �猌����R��!@����u�Ŝ�#b*"���G}��K.�T���Ӟ�xL4�?)�D*�?��QOE ����?_;  `��dǎo9p��skw   ��bii�v '�hD|$�4�R����ۏe�}��߻�>�&%Q4c��qp�ئ��
��(�(��b ��e��/`������f��""8�dl<�������:���U��>����n5)�ه�z��y��ݬ�&?l@w��z�����?� ��>��VJߊ��v�G���n���>>�յ��   �	�   ̤N�c�0�^��o7M��ib0�F�_ǃ�06��@���K���FD|���7M����T ��&"v��rg   ,$w   fRJ):�N�F��) ��ߎ������`���>�v���������u pI�}����^���4ߎ��v��V�����;::�����   i�O�x�w�rgg�Osw   ����I4M�;��3���'"�*"��K/����~��'�� ���[������_�i��.|�	 �������`  �Kb�  �L��QUU� ��4"�>"~�R�q����{�����Q �Y�Oh����o��oG������˵��[�۹3   ��;   3���4�Ν@ӈ�ED�8��A���O�q�;
��t>h��T��L�[�j�. ��t:������t:͝  ��Z�   ��t:���3 ȣ��7#�ͦi���hT��������n����o��M`Q��G?j5M��#��G]����M�4 2���3n  �d�   ̼V�EQ8����""�������8��N<8��'M�|�����?��?��`���?�R�?)��&�o�������l��qp�V�  ���r|�w�y�/wvv�4w   yM��8;;˝�|��_�r����`p�;
�������S�ߌ���&�M��҃�� �Wܸy3�n�Ν  ���  �\(�2Z�VL&��) ̾�#��ͦi""�����aD��(��|����YD4�b?�яZM���T��L����������98
�lΆC�v  �+b�  ���v�� <�2"�<��C]�1�"�o#�oSJ�4���[Y+�P��{�3-���H��6�H��[�y�}O9�,6��r'   ,w   �FJ�)� \�ߊ�?��?yxr�`0؉���R��i������ <����_jE�A��V<������������ݿw��˝  �4�  �+�n7��i<#�z=~u��?9���/~���|�;g9#��{��R�(�)��4�[EJo5�)w �i���   W��  ���R�N�UU�N`9�o4M�""�޽;��oJ��SJ�������wO�f,���ݕV�RJTG�Q*�?�����(#�?��+ �i�֭8;�+  �U2p  `�����Q�u� �O'"�_o�&������;�aD|�R���j���o���7`���?��J���"��RěM�|5R�zDt�8?��'9p���i�����   X:�   ̥n���, f���'�'M��x<��`p;"~����(>������������NY��D����W���j"~?��#"R�� [;;1�Lrg   ,w   �RY��j��d`�}9"�y~=��{���#�SJ?��l�槃�����Bz��w;����狀���4E��4_k"^m�OcO)�s��5��0n��   XJ�   ̭N�c����BD|#"��p�1�#�zD�,��a�4?m���������	�L~������?m��Շ����ތ�uݍ�'�7�1; sa}s3�ov   �����;��;;;��  ��TUU���� pYv"�ϯ���~4��VK�����J�(ތ����7���jJ�kMD?w \���Ǳ���;  `i9�  ����vc2�8Q�E�������`0�����RJ?M)�����?��w�s��X0��n��W_��E��^�����F�W#�͈x���k""Rr*; ������Ν  ���  �{�N'��ʝ W�����M�D�4q����`0X���{J�gM��4"V���T�������������N��Rz3"�H_m"~7"�H3�a� p�v��c4��   Xj�   ̽V���8�Ν ��"����p2�#�Z�r���EQ�N�Ӎ�`0��\����_�D�Q��?DJ����璉~/"�Ť���"��!�'a XV��(���sg   ,=w   �^J)z�^����N�Y�JD|��z4~�N��>���k]������{x{�4o4o���o4o<z�i"9� >��֖   f��;   �(�h��1�s� �<�̓����x0~߈���XO)m4M��w��%\�>��7ʺ��&�7RQ<�ǃ�?�TU'�/O_��+ �d�����Ν�   ��;   ����t:u� \�Wϯ�?�������`0���`��Rڎ_��3��2�ɻ��y��W���i������N`�JD��<"�E)��)��z#v x1u]���V�   ��  �P��n����� �eӎ#��#⭈�<~���~��ה�NJi���p<���{���W����&�+M��"�i<�~������H���� Khs{ۧ  �w   JY��j�b2��N >���B�4��_���؊����L)�7M�����a������߬����������JD��4�WRJ��c�/G��?��~�� ����4n�ʝ  �c�  X8�n�� �W7~y�uD����O8?�����aD�G����oEĭ�(�>�v�w����ݾ�|�Տ��/���ߊ��H���Z�4��"�ID�FD�������WF|����`��� �}M����F�   >��  ���R�n�UU�N .W�y~�Zu���쪪b0DD�_w>����)�G_K)������ID�������I?��_������R��+��+Mė"╨�W��x5���T����ă��k����8�;q ���A�����   �Sf��e�y睿������   ̟����N��3 ��tv~��#�����_��aD�FD����5MsQŽ��DĤ��{�v��(�QUU�"�������}vv��p8�BY�+�rQ�_��z�r�4_��V"��4_�S�B��+)�W���z����r��  �c4�O��GC  0;��  ���v�qzz�; XL+�׫������Yê�x����'�����7������_h����7���;M&)��'�}�(���}��(SD;Rz9""=����#"��BJ��C|������������{�ǭ��VJ�̓����G_OM���_�� x:[[��   3��  ��UE���O��  �˟�����O���8���QO�E)���?���<6:������1J r�}|�w�|�O   �'�)6   ̹n��猸    X��$�77sg   ���  ��z�^�    f���fL&��   <��;   �(��t:�3    ����q�>>Ν  ��0p  `)t:�(
o�   ��d2�����   <w�  X�^/w    �on�d2ɝ  �S0p  `iE�v;w    W���q�>>Ν  �S2p  `�t��(
o�   ��d2�����   <w�  X:�^/w    W`}s3&�I�   ���;   K�(�h�۹3    �D������q�   ���;   K���FQx[   ����q�ol��   �9��  ����z�    �776b2���   �9�  �����N��;   ��pw��͝  �s2p  `�u:�(�2w    `8���N�   ^��;   K����N    �5M�7oF]׹S   x�   ,��R�����    �lmo���Y�   ^��;   DDY��j�rg    ��޻{�3   � �   p���EQx�   0O&�I�\_ϝ  �q�   ��vs'    ��77c4��   ���  �cʲ�N��;   ��p��0n��   ��  ��t:�(�2w    O0cck+w   ��   >C�׋�R�    >C]�q}m-�Ν  �3p  �ϐR�^��;   �ϰ����0w   ���   ~��,�����    �1�GGqxt�;  �Kb�   O��t�,��    D�p8�����   \"w   ��^/RJ�3    �Z]�q}m-�Ν  �%2p  �ϑR�^��;   `���؈�p�;  �Kf�   O�,��t:�3    ����aݾ�;  �+`�   O���DY��3    ���p�[[�3   �"�   �z�^��rg    ,��t�kkQ�u�   ���;   <��R�z��    K���F���   \!w   xFeYF��͝   ��vvw���q�   ���;   <�v��v;w   �B�{�^l����    w   xN�n7��[k   ��4��X][˝  @&��  �XYY��R�   ��P�u\�q#��i�   21p  ��R�^��;   `!����p8̝  @F�   ��ʲ�n��;   `���������   df�   ��nG��ʝ   0��޽�;;�3   ��   pAz�^�e�;   `��*Vo�̝  ��0p  ����"��;   `.L�Ӹ����4w
   3��   .PJ)VVVrg    ̅7oư�rg   0C�  ��Ea�   �9�77��ݻ�3   �1�   p	ʲ�n��;   `&����[�3   �A�   pI��v����    3��{����;  �e�   ����FY��3    f�p8�յ�h�&w
   3��   .Y�׋�R�   ��&�I\�q#��i�   f��;   \��R����    ��u�o܈��r�   0��  �
��bee%w   @776���I�   态;   \��,�����    �Rۻ�qt�v�   愁;   \�v��N'w   ���ux;���3   �#�   p�:�N����    ���ݻ����;  �9c�   t��h�Z�3    .���i���E�4�S   �3�   �I�׋�,sg    \������j�u�;  �9d�   �z�H)��    ���4����d2ɝ  ��2p  ��RJ�����  ��W�u\�~=�U�;  �9f�   ���bee��   �[M���7���4w
   s��   f@Q���rg    <���͸{�^�   ��;   ̈�,��  ������sg   � �  `��Z��v��3    ����A�����   `��  ��i����trg    <���Qllm��   `��  ��t:F�   ��:�s'���sg   ���  `F���h�Z�3    >��ݻ����;  �e�   3*��^��   �'''q}m-��ɝ  ��2p  �����,��   ��;=;��WW����)   ,0w   �+++F�   @6UU��ׯ�t:͝  ��3p  �9�$w    ��h]���$w
   K��   �DJ)z�^���   ���F�k�b4�N  `I�#   s$�+++F�   ���L&������   \)w�  `��   �m2��/�]�aU�N  `ɸ   s��   �,����a�   ����   0���  ��f�  f���    IDAT@n�  �{8rO)�N   ��d:����  ���   �\J)����;   ��&�i|���qf�  @f�   � �܋�[}   ��L&����u�v   f���   � RJ����$w   �M���xu5NOOs�   @D�  �By8rw�;   �y&�i|t�q;   3��n   X0EQ8�   x��d}�q����N  �O0p  ��R�~��$w   �W�F������p�;   ~���   ����˲̝   ̈�h��v-�U�;   >��;   ,���'�   1����(w
   �Z�n  �p�;   ,��p]���8w
   <��;   ,���#w   XB����k�b<��N  ��e�   Kdee%Z�V�   ���?9�_\��v   愁;   ,�^�g�   K���I\[]���s�   �S3p  �%�����n��    .���������N��S   ��8�   �T�ۍ�(����)   �:<:���4M�   xf�   ����n�   �awo/�vvrg   �s3p  �%�n�#���0w
   �6��co?w   ��"w    �_�Պ����   �sh�&nnl�  ��  ���(�2��~��r�    O���~�F�:<̝   ��   x�(�XYY1r  �90�L�����ݻ�S   ���   �PE���(
l    �j<�G׮���I�   �P�T   �"��~?ʲ̝   |�p8���Q���S   ���   ����J�Z��   ��{����?�8F�q�   ��P   O��v�(��F�S   `��>>������:w
   \w   ��RJ��t�(���s   �b�� 6��rg   ��3p   �J�Պ���8;;˝   K�i�X�܌[���S   �J�   ��Q�e���H)�N  ��W�u\�qø  ��b�   <��(bee%��+   �e���?�;w��N  �+�N4   �̊��~�eY�N  ��s6��?�(N��r�   ��k�    ����JTU��8w
   ,�������ZL���)   ���;   �B:�NEUU�N  ��v��0�77�i��)   ���;   �BRJ�n��(��n�  �3j�&6��c�� w
   dg�   \��,cee%��a�u�;   ��d2�յ��w�~�   �	�   ��)����}:���  ��v6���ըF��)   03�  ��Rz4r�L&�s   `&ݹ{7nܼ�q   �w   �R�z���QUU�   �)�����;   f��;   pi��v��b8�N  �욦��qxt�;   f��;   p�Z�V���8;;��ir�   @��$�������s�   �L3p   .]Q��K/���YL���9   p�NNNb����F�S   `��   W����d2���r�   ��8�};nnlD]׹S   `.�   W&��v;�������9   pi������88<̝   s��   �reYF�ߏ�p�;   �x<��7n���i�   �;�   @EQ<�O&��9   p!�߿�7o�x<Ν   s��   Ȫ��FY�QUU�   x!�c}s3��ɝ   s��   �*��v;����ph   �ܩ�:�77���(w
   �=w   `&�e�~?��΢���9   �T����7n��p�;   ��;   03RJ�������ǹs   ����܉����N��S   `a�   3���FQ1��i��9   �	M����n����N  ��c�   ̤v��V+��΢���9   ��8V�����$w
   ,$w   `f�����GUU1�s�   ���܉����N��S   `a�   3���FY�1s�   �����������͝   ��   ��V+��~�è�:w   Kb4Ǎ���r�;   ���;   07��x4r�L&�s   Xpw�ލ7o�t:͝   K��   �;�^/&�I���)   ,��ibgo/vvws�   ��1p   �R��zt�{]׹s   X��(Voތ����)   ���  ��UE�����*��q�   ����㸹���4w
   ,-w   `�u��h�Z1�i��9   ̙��c}s3��r�   ��3p   BY��Ns�L&�s   �����z�fTU�;   w   `������FY��	   <Q������   `��   %��v;ʲ��pu]�N  `ƌ��q�fܿ?w
   �)�   �B*�"��~TU��8w   3��ΝX[_��t�;   ��   �B�v�Q�eTU�#�  ��t:����8<:ʝ   <��;   ��Z�V�e���	}   K���$���cXU�S   ��a�   ,��R����d2q�;  ����:v��bwo/w
   ��  ���4w  ��pvv7�����,w
   ��  ���R�^���$F����  H�4���ۻ���  �2p   �RJ)��v�eUU9�  `�øq�f�:�   斁;   �Ԋ�������QUU�   �ӭ����ڊ��s�    /��    ��i����  `��F�X[_�{���N   .��;   ���(����h4��h�;  �'h"��֭�����2   ,w   �O�t:�j���  0�����Nm  �d�   ���>�����9   DD�4Nm���@2   ,(w   �'h�ۏNs�N��s   ���p7�����4w
   p��   >GJ)z�^L&��  \��ibo?�ww�i��9   �%3p   x
)%��  \����X[_��p�;   �"�    � �+++1�L,   .I]ױ���{{�S   �+f�   �Z�V���KQUUL&��9   ��{qsc#F�Q�    w   ��R�^���4�����s'  ̭�d���qxt�;   ���   ��e�~?F��  ����۱����    w   ����t��jEUU1�Ns�   ̼��0nnl���I�   `F�   \��(����t:����i��I   3�����ߏݽ=�   �O0p   �`)�h�ZQ�e�F��ǹ�   fƝ�wc}s3F�Q�   `�   \��Rt��h�ZQUU�u�;	   ��d[��qxt�;   �a�    ��,����1��P  ,��i��֭�����/   ��   �H�Ӊv�UU�d2ɝ  p��߿�[[qvv�;   ��    W(��^/��iTU��B  `!�����ىã��)   ��1p   Ƞ,����1�����9   �i�8�u+�vv<�   <w   ����v�Z��F1�s�   <�{�����V���)   �3p   �,��n7Z�VTU�C  `��F���ݍã��)   �0p   �eYF�ߏ�xUU��  x���c�� v��<�   \w   ��n���j�h4��x�;  �W߹[[1�r�    ��   `�����F�ݎ�h��$w  @������V�?9ɝ   ,(w   �VE�z��N�QUU�u�;	  XB��8�ww���a�   `��   ́�,����x<��hM��N  �@]ױp���1�Ns�    K��   `����h��QUU����9  ��}|���1�r�    K��   `u���t:QUUL&��9  �99=����89=͝   ,!w   �9�R�^���4�����s'  slXU������s�    K��   `Εe�~?&�ITUM��N  ��d:����8�u��	    ;w   ��j���j�x<��hd�  <Q]ױp���1�Ns�    D��;   ��i���j���  �i���(�wwc<��   �w   ��Rz4t�FF+  @DD�>>����   3��   `������F�Ӊ��b2��N  2�{�^l�����i�   �'2p   X)���zQ�uTU��4w  pN��bsk+�ݿ�;   ��   ,��(bee%��iTUu]�N  .���b{g'n�N   x&�    K�,�GC��hd�  b4���^E�4�s    ���;   ��J)E�ՊV���$��2� �95�b�� n����   �\3p   ��  ��d:�����?8��L   �B0p   �Cw  ���$��  ��c�   ��x8t��1�� `FL���;8���}�v   `!�   �k���h�ۆ�  ��t:��[�bw?��i�   �Kc�   ��z8t�F1�� ��<<�}����   X
�    <�N��N'&�ITUe�  �d2����[��   ��1p   ���Z�h�Z����ػ���&�yцP���/�5�E�D����)�VC�pN(�����I ���m�����   ��	�   �n�C���8  �꺎?��b�\�s5   ���    ��ס{�4�u�Г  �&��:>==��b�;#   ��   ����w]u]� �+N�S���S<���   ^�   �Ӎ����߄�  ��~���?}��z=�   ���    |�K���}4MM�=	  �����?���f3�   ���    |��h��<�ө� ��QJ���*~��8�NC�   �	w    ~�K�>�͢mۨ�:J)C� �����X,��ǧOQ{s'   �7�   ��UU��4���5t��~�Y  �Cڶ�O�E<-Ѷ��s    n��   �AM&��L&Bw  n��|�O�E,�K�   �Aw    R���]�E]��u�Г  �m����X�j�z
   ���   ��x<��~�-J)Q�u�m���g @DD�R�e���?}���8�   ��#p    ���b>��|>��i��k�;  �i�6�e|Z,�i���    �-�;    �M�ӘN�Ѷm4M]�=	 �q8�i��痗��~�9    wO�   �͘L&1�L���h���L  >D���zO�El�ۡ�    <�;    7g4�|>��lv�K)C� ��u]�������z   �C�   p�����l��,ڶ��i�뺡g pcN�s<-�X.�����    <4�;    wa2��d2���i�h��Uw  �����:�el�ۡ�    ��   ��2�b>��|>��i�iW8 �j�&���xzz��w�   HG�   �ݚN�1�N�Wݛ�z  (��nc�\�j���~    �   p�.W�g�Y�mu]��  @�u�|~�?������    �/�   xUU]���m{}  p_v�]<}������s    �w    �d2��d�W� �@۶�Z����SO���    ��    <��Wݻ���i\u �%"��m,>_k��E   ��'p   ����q��㈈h�&�����^ �[M����9�e��z�9    �Dw    x��{���� �am\k   �{w    ���(��y�f�h��Uw �_�t>�r����s�m;�    >��    �������~��] �������*��ϱ�   �/$p   �o4�b6��l6���i�h�f�Y  7o���b���z퍄    J�    ?`4�|>��l]�E�4�u�г  n��t���K,��h�v�9    L�    ?AUU1�Lb2�D)%ڶ��i����� ��4M��V�|~���8�    �   �OVUUL�ӘL&���5v xd}��j����sl�ۡ�    ���    >HUU1�c<�|>��m��h�6J)C� �p��Xo6�Z��e���m    ���    ��L&��L&����  �'%"��}��V���m�=	   �"p   �\b�RJt]M�D'� n��t���K,��h��   ��$p   �UU�E�~��.v n��t���*^^^�t>=   �; p   �$����t��4J)�4M�m}�= ��|>��j�//q<���   ���   @BUU�l6��l}�G�u.� ���:V�u��V��   ��   @r��(F����{۶bw �ÝN�x^��e���K�    �"w    �!UU�t:� B�   ���    p����]�E�4bw ��\����8��C�   ��	�   �TU��$&��5v�\w x����.V�u���h�f�I    p%p   �;�:v��/b�R��� �!t]��6֛M��V���Г    �]w    �s��8��q�������� ��u��6V�ul�[ot   �&�   ���F���f1�͢���u��놞 ���)�W�Xo6q8��    �L�    j4�h4��t��/bw^�6�}��66�M�6�h�f�I    �C�    @TU��$&�?���uw ȫ���l��Z�c��zc    wE�    ��{��/��� ~���c���z���zu]=	    >��    �G�����s���p�   �G%p    ��{��/��� �O�u��n�W�   xTw    ໽����� �WJ�����6��]lw;��   ��    ?������ ��꺾^h_o6���Г     �;    �a^凜������ �wM��n���M�=	    ��    �DUU1�c<GDD)%ڶ�F凜���i�6��]l����vq:���    7G�    ����N�1�ϣ�]�].���%h�������p8=	    n��    H����L&1���ז�w �i�6v�v    �Pw     %�; Ck�&v�}l�����q:���    wO�    ܄��}�G۶�w ~H)%��c��������n��g   ���    7��GD�f�������+凜!'�X�u�?b�����s�uC�   ��'p    ��h4��h��4"���~y���꺎�~�E�    �#p    �������{DD۶��}�}m�����u]��/����    �A�    <�ױ{�_W����^z�v�R�|>�n��^h?�NC�    ���    xh�+�].�����t:��x�����!��C�R��    �$w    �7F�Q�F�/����{��.x��9�ßA�~����_    �sw    �������{���|�RJ���/.���   �1	�    ��{��K)��.z�K�uq<����t����k%    w    �����/���?�����ܳRJ��:��#�����!�z    ���    ��UU��8��qL�������_�w�[�4MO�8�N�����k    ���     �F1����%|� Z۶q:��p8�   �!p    H�k�{�u�k��wࣔR�\�q<�|>ǹ���ٻ�z    p��     7b<���{���5��i�6꺎��������(�=    xPw    �WUU���𥔯���Uxm�ƹ����8�O�s��g��   ���     w�����*F�ѻ}��폁�PJ��i�t>���/�"v    ���    �%|{�="��_?�F���i�\��|~���k�^7��&   ��"p    �o����x�n�~�O������m�/���i�?���wU     ��    ��2��W���:v/��s�JD�m��`�m�k�~yn�&��z*    @*w     >�?�ﯽ��/ת��dTJ��m�뺨/�z]G�*f�\a��-    ���    0�o�#��k�]y�7�����z�F����h���ǫ�     �8w     n¿�/���o��~���m��>�������k���F��    ���    ��TUUTU�]��:vȿ�񷯽}�/�}}t��ϱy)���W�F�o����     �w     x�G����R����^�/������|)忖��_��J�(    IDAT���w�>�u�u��s�����y�Z�uїQJ�����    �{�     ��.����E����������    ��=            "�           $!p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          H!}�~>�z           /}�����?Co           ���          xw           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���      �v�ئa( �hl��PDM����؆	�Af���'��7�   @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	���l���,��������y����    p��<=\.��;    �?������>���it�=뺾L��:�          �cͣ           �t2�          ap           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��  ���    IDAT        @��          ��;           	w           ��ˮ�0<�%P���*B^��1�`,          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          ��9pg������           ����Z����           �Y��           0cp           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p��];&B �0��-�w��o�s�U         �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��        �WA�    IDAT  ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @�m:�g����   ���t    ��.�   �����~�s��           |�u:            �2�          ap           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��  ���Ko�i��|���)Mg�fQ$���ŰDH���lA,��8H0�,1����q�ĉO,`�X��j�����>�mE������       �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "Z  X����z��z���a�W���e�ޢ�7�n=�{q3������;{�[��>s���~}s��z�x|U��e� |�<�U����������;�^����� ��� �N9��N.Z�`ÞOj��������NZ�`��p~O�������㷭g �ٗ���xr��N���3 ��z}T3�$����uN����� hJ          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�     �揓{5[������m�[u6��'��gl�_����l��X��E���8i=X��������-���y�[5t�\UϦ�lz�z��n��� ���    ��\�����F7������u2����U/n����
X�ٲW�>l=���U=>�n=��̆ާ  �w�k=            ��           ��          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          a�z  �:}uuTϦ�gl���I��nZ�ت=xU��k=���ZOغ����������.��'   �w����ً�3`�~��~�φ�g ��O�����X�7�a�����3 �� ;�f٫�e�~�f�������\�5��^]���  �����d0k=�n����0�/�7�sn�� ��^          @$�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �       4�j=    �1h=      �g>o=�����������φ�˗g�g  ���ZOغ�=z^����  v��          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          ���  x7W�~Mf��3��x8�^�Z�`�����w������z �_&�AU��E�:�[�`��{˺7����UW�~�V��a���V��_�]5�;u�s���]��-�p�h=c�F��}��^��. �D�� ����>o=b�~��u����|X�z��� ��~��;u���h�޲>��Y�l���U=_���U�}�A��z�z���`^?~���`~���5[v��Y��/�Z�ت�����Z�ت�/�����3  ���cK           � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p        ��k�6� EA(�]6c-�C�6$B�OX��/p��pa� H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          �p3{   |��q;��������@��t;����g���r5{Zƕs͟�~�̞��^?����̞�,��X�qٸg�қ `��/�n�{:��w           ����           `�; �H�    IDAT          w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	���|>ogo           `}��}��0{            ���;           ���          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w          �d�nw�H���������ﯕخ�z�mv�N�!�ry	%!к��A��VA�          �*�          X�;           � p          `�           ���          �U�          �
w           V�L=���y~*��>vY�o~���           �����i�_��͡����C����|Ώ>          ������-eY�ͯo�����G          p�y���4M��yY��
��C�e��e��2����)_�          `M.��%P�կ�%pO ˲(��_?����g�          xK�4}����͟�$\�]��\������}�>M�?.�          \|�_~���l��W��k�UU���������          l�<�1��������J�a���M�u�����          �z]��K�>�7!�5�߰���������_^~@�          i,��M���e�������y���K�~	ޅ�          ��/WٗeI=�C��m�
߿��>M��          ~����}߿����
��kY�EQQ���.���o�4%\	          i,�}��0�\f�E��M���;          [t	���	��=w>T���y���ӻ\z����4Ų,�W         �������0�a�����~t������          �-����}]��<ϩgm�����>z�>x���O�          ��iz��]g�wV�GW�/��<�1��
          ��%h�.���qSO�9w�R���yDD4M�<���;          ���A{�u1MS�I7O��&\������_���4��         @L����}/h_!�;�t	ޫ���;         �-Z����0��Ŀ�s��/��8�1�s�u          ��eYb�o��s]�ܤ�(�(���:�e�&xw�         �z��]�E۶�u���WN���˲,ʲ��,�i���9�q�i�b�g�;         ���m�F۶1C�9�!�;|'���:"���%x�         |�y�_.��Ҿmw�����GDL���{`         x?�4�\i�.�>��^�(�(�"꺎y�_.�OӔz         ���!ڶ����8��Cw�Cy�G]��,�K���         ��,�]׽\j��9�$��Ȳ,�����bY���}��X�%�<         ����+wxcY�EY�Q��������(v         n��Q��|�T�SwxgEQDQQ��7�;         ��-���w]'j���|�}��!�iJ�         ��t]��٥v������˲�4Mbw         �j�}����zWL��}}�}Y�����        �5��%jw䗷"p�ɲ,�����b�����s          k0�s�m��1�aH=���J�yu]G]�1M�K�         �e����|>G۶���p����(����}��Գ         ���>N�S�m�[����dYUUEUU1��K��'�         ��0�s�m��1�aH=�$p�+��y�u��U�i�R�         �P�uq>��|>;�KRw؀�,�,�X�%�a�q�         �K�4��|�����.�!p�ɲ���4M/�;         �E۶q:��m��S��QEQDQ1�s���0x�         �Q�<��|���g��Y5�;l\��/W�/��'&         ��0��x����P.WA�7�,�(�2�y�ab�ԓ         �7�,K���8�ZA���nP���4M4M}��0~*         ��<�q<�x<�<ϩ���Í��:꺎i������)�$         ��a�������[�������(b���4M1���$        ��k�6��ct]�z
��;���(�(���:�a���SO         ��<�q:��x<�4M�����?�eY�uUU�01��-        �D�y�����1�yN=ލ���K�^�u���0��/         � �8��x����P-7A����,�,˘�)���        �;��%l�["p^�(����1�s�}�8��         �жm<??G����@w���y��.�y�abG/         �m�xzz�aRO����_��<�����bO�         ���-�;�f��         ��ey	��qL=VE���K�^�u�}/t        ��o�~:����9�iJ=VI���,˄�         ����v�w��}���˲��         �N��#p>�%t��*�a�        �Ym����SÐz
\�;���<	�/�        `���w�@2y��n��i������)�$         �#}����c�}�z
\5�;�\Q����         \�q���)��s�)�	w`5.��8��u],˒z         ��4M�����)���;�:eYFY�1C�}/t        `5�y����8��6xw`����&t        �T�e������1�s�9�Yw`ղ,��������>�aH=	        ��u]��1��<�;p�,��i�,���>�iJ=	        ���1�Ct]�z
��;pU����~�8F��^�        �77�s<==��xL=n���JeY�\s��>�         6`Y�8����˲��7I�\��������>�aH=        �+�u]��1��iw��eYM�DY��u]��z         Wb��xzz���z
w`C�������k�^        ��Y�%������Yo+"p6��먪�%t        ���m��!�iJ=���ؤ,ˢi�(�2���y�SO         �i��p8D۶�� ?!p6�(����������s         H�x<���c,˒z
�w�&�uUUE۶^R        ���1C�)�o�7#˲���1�ct]��         6l��xzz���z
�
w��eEQD�u1�c�9         ������!�yN=x%�;p��,��n�4E�u��        ؀y��p8��|N=�Cw�Ewww��}�}�z         ��v��;@D�uEQ��        pe�i���mۦ���;��r�        ຜN�8�,K�)��|�5w        �u��)���S�7&p���        ��|>��pp�6J���k�m�z	        ���y����h�6��	��EQ�?��?�u]Ðz        ��i�6\m� p�MM�DY���        |�y��p8��|N=� w�W�\so�6�qL=        `���������)��	���n��q��:��        ����S<==��$ p�CeYF��Ѷm��z        �՛�)������S�D� !�󸻻���}A        ���sG��	��@]ב�y�}�+        �W��9�C����S�����,�(��.�qL=        `��a���{��B����,��n}�G����         ���t���˲�������uEQD۶��        ��Gw]    IDAT�,�����9�`�� �(������mc���s         ��!���c��S�����,�b��G����}�9         ɜ��xxx�eYROVL��꺎<ϣ�:_�        7eY�xxx����z
p� �,�(�"ڶ�i�R�        xw�8���}Ðz
p%�� nI�e����S         �U۶���'q;�*.�$�4M�y]ץ�        �枟����1��
	���*�<��mcY��s         �ڲ,qmۦ�\�<� �[VE���E�{8        ��8����G��E%@bY����]���         �S�u��ӧ�1���	�Vb��E]שg         ���x�ϟ?�<ϩ� �\0���uy�{�        `��e�����)�`C\pX��,���.��C4        �N�<��ϟ����SO�P����(��S         �1C��?����SO6H��RY��~���,SO        ���������1MS�)�F	�Vn��E]שg         7�t:ŗ/_b���S�s�
�uY�E�u��         7���)���R� n���JTUy�G۶�,K�9        �X�%�|>��܈<�  ~_Q���#˲�S        ����9>�,n>�����ywww���       ��1MS|��)��O=�1�H�+�eY���(�"�        `c�q�O�>�8��� 7H�p��,��neY��        l�0��ӧ��)��F	����        x+]�ŧO�b���S�&p؀�nUU��        \��m�˗/�,K�)��s�`#���<ϣ��S        �+r<�p8��w�M�\q�        ����9S� x�� �۪�*��I=        X9q;�F.�lPUU�eYt]˲��        ����c<??���.�lTY�.�        �p8���j	�6�,�����g         +�����1����l\Q"w         ����t:���Kw� r       ��v��9��%p�EQ�n�K=        �`�v�j�nHY�"w        �!q:�R� �mw�#r       ��p8������ �;        l��p���z��	�n�%rϲ,�        �=>>�ہ�%p�aeYF�4�g         o���1���S� �cw�'r       �m8��v��	��������3        �?t:��p8����� DDD]�QUU�        �+�m�g �	�; /���       �i�6���S� x3w ��4M�e�z        �/������X�%��7#p�v�]E�z        ��8Ɨ/_��������ny�i        �f�����s��z
��S.�CY���       `e�e�/_��4M�� ��" ?��y�v��3        ����}��S ލ��_�       �:<<<D�u�g �+�; ��,�h�&�        �YOOOq>�S� xww ~KUUQUU�        ps��s<==���!� ���i�,��3        �f�}�g |�; ��4M乧        xo�4ŗ/_bY��S >�B�Wɲ,��}dY�z
        lֲ,��˗��9��%p��.�;        �>�|��0����� ��<�c�ۥ�        ����]ץ�����?V�e�u�z        l��|�����3 ���W꺎�(R�        ��7C<<<����������"�=�        ����9�|�˲�������eY�v��3        �j����4M�g $'p�M�yMӤ�        W���1��K=`� �����,��3        �j�m��ϩg ����7���"�=�        ����)R� X" on�ߧ�         ��,K|��%�yN=`U� ��,�b�ۥ�        �����0���:w �EY�QUU�        �:��9��c� �$p��4My�        .�q�����3 VKu������eY�        �ܲ,q˲���Zw �U�e�4M�        ����SÐz��	�xweYFY��g        @2}����s� �'p�C�v��sO;        ܞy����>����4��4M�z        |����4��p� |��(����3        �ÜN�8�ϩg \�; ����sO?        l�4Mq8R� �*
C >�n�K=        ����},˒z�U����<��iR�        �ws<����3 ����$ʲ��(R�        �77MS<>>��p�� $�e�+�        l���},˒z�U��L��"w        6�x<F���g \-�; I�eEQ��        m�x||L=�	�H*�2W�       ؄��˲��p�� $��yTU�z        ����]ץ�p�� �B�4�瞖        �>�<��pH=`�� �F]ש'        ��=>>�<ϩg l����(�2ʲL=        ~[��q:�R� ��; ��4M�	        �[�e�����3 6E���dY&r       �*���1��M��:UUE�{�       `��i�����3 6G=�*��       ��=>>Ʋ,�g l���U*�"ʲL=        ����8�ϩg l����r�       �5:�' l����ʲ,�N=        ^���!�����ju]G�{�        �y����)��MS�zUU��         ����<���iw V��*W�       Hj��8��g l�Z��P�u�	        ܰ���X�%����pʲ��(R�        ����9��� p�j4M�z        7���1���!p�j�yeY��       ��.��K=�f��*u]��        �q��c	��*y�GUU�g        pڶ�aR� �)w ��+�        |����� n�����eY�e�z        v>�]oH@��Uj�&�        6���9���$p�*eYUU��       ��������U�u�	        l��� ���Z��       ��\oHK��U��*�,K=       ��p� -�; W-��(�"�        6��:���p��N=       �p� =�; W�w        ��0�u]� 7O��&��       ��p�`� lBQ��       �G�i����z !p`CʲL=       �+�z;�z�،��"˲�3        �"˲���"w 6����        �"��)�yN=��%p`S�        ���xL=���ؔ,ˢ,��3        �]��8��g ��; ��;        ���v����9EQDQ�g        �b�4E۶�g ��; �T�e�	        ���� �$p`��        ���|N=���IY���       ���mc���3 ��; �UUU�	        ���tJ=����YEQD�{�       ����]ץ��O�� ش�,SO        `EN�S,˒z ?!p`Ӫ��,�R�        `%N�S�	 ����M˲,��H=       ���>�qL=�_��yu]��        �
Ðz �B����v�Ȳ,�        Ӑ ����ͫ�:��I=       ���y��(D� +'p`�ʲ�,�b�ߧ�       @B�<G�e���RO�� lZUU�4���       �Q˲Ĳ,�ߎ����Yy�GY�~�       ��}��e�Ҕ �>w 6��oD��}�%        �4��7v(`�� lVUU���i��sO}        ��r���i�Ȳ,� ~E��&E�Ø�i�k        He���Y�E]׉�+w 6�����1       �-�<����� �;� lN�eQ���n���        R�Y�^U�O ���9u]G�e?�;//       p;�e��߻��>w 6��~��7&        ��g��/����!E ���)eYF����i�Z       @J�v�=�2�VF���TU��S�eE�k        HeY������?` �K��fEeY��Ǻ�       �m�v��"������ �� l��\o��       l��\o�p�`=� lB��}�="��-       �������V|M{����	UUE�e���^Z
       `��eyU�qww�Nk x�; W/˲���՟�4�;�        �y�_�9u]GQ����p�^{���w       �mz�����~��K x-�; W�OC����(�       `��4po�&�\Z	��Ga �ڟ^o���       ؎eY�8pϲ�w��� \��i������;        �4��_}�n�s� !�� \����!p       ؚ?��~�eY�v�7Z�k	��JY��I�^��_G�        �������w�D<�p�ʲ|�o"�,��(�`        �-��&�{�e����` �%p��������g       ��[�����w�<�pu��z���  �?{w��ƕ��v���A�F��+���l[,����6�eY�:+#Ba���xmS �`     ��[�!p`v�:Ho��M?        u���w������m���4�R"���       ��K)�j��=��������c���i�7��        ��8�1����b��7�� |��������.��m�.       ��x����+� �#p`RJ���       ��=���i�w�� ��; ��uݻ]o��        ��{����]?> �%p`�r���7M�=        �k�w��m�:�pw &����<Nξ,       �m���?% �VJ��iN�Xm۞�q        x[�8��qJ)�\.O�X �J��d��b�X���N�       �a8�c�V��Y~	�^<�0Ym۞���R��       ��s���=ڸZ�N�x �F��$���뺓>f۶'}<        �i�XD�4�g �%�; ��u]��N����        ��S^p�^�O�� �@���RN~�=�W�s��       `nj�m�F��'\�s��`rj��w�       `^j��/��u���=>�9�0)m�F)����|l        ~^��=�������#�; ��s��bQu��       `^j���"�����������jO�       �Ӯ��jO 8w &�i�h۶��       ��ajO��ib�\֞p� T�R���kψ�       �5��J{�� T�u]�<�/I��        ��qkO���y\�׵g ��4jB .V)%���=�o��       0/]��b��=`�| T5��w       �y����ϭ�k�	�o�
@5}�O���7       0)�����=`�| TQJ���j���RJ�	        �X۶�X,j� �%�; UL���        �0C�	ߴ^�u( ��3' '����_�Oy        �R�����3 fG��I�R�m��3�U)��        �@�u�X,j� ��; '�R��r)��S����       �_�8֞�]��:���=`6� ��b��E<��/�        ���R\__Ϣ�� '�4�w�       ��p�="���ժ��Y���rα\.k��a.�       �֖�e�m[{��)� xw�Ţ���"p       �=\__GJ���IS�𮺮�RJ�?�7        ���s\__מ0iw �M)%���=㧥�D�        ����b�\֞0Yw �E�9���lC��       `���u�m[{�$	�x}��:Ǳ�        �c΍���u�,���gF �\���4M��e�q>        ӗs�����3 &G���*���I        �����rY{���x3)�X,gq���        ���z�$�g� ���r9��       ��Ǳ��7sss���3 &A���X,g�"�w       �i;��#����g���� ���m��$        N�.�GD4MWWW�g T'pුRb�XԞ��       `�α����,[��!p����b�\֞�.���        ��\�����h۶��j� ������	       ���s�r}}9K<�����_�X,��R{ƻ9�w�       0}9總�=��[� ����i��3        �l�R���������S�����k�xw.�       P[�u�^�k� 8)�; ?,��Ţ�        ���R�\�; ?$���2RJ�����        L���U�m[{�I����R�V���r�l�       ��R�5FD���D)���ww9�" �l�X\T�>C�	        �7)��������L�� �W��"���=�\o       ��K���s���ۋ��.���o��>ڶ�=��\p       `�J)qss#rΖ���j�6���=�
�       ���m�����w!p�����bQ{F5w        ����X�׵g �9�; SJ��="b��        ໖�e,���3 ޔ��W��X.��R�=�*�;       �<�,�\���8/�������_,�G�       ����������7!p rα\.������        �\__G�u�g �6%#��K)�ۿ0�c�	        ���R�	�r}}m�֞�[Ԍ L��u.�       0G)������ijO�e�F����RjO��;       �<���O"w`�� H���a�=       �$r������-�;�����        ����]'̍��¬V+/Z����        ��������V/̊������}�á�        ~���߉܁��\��R�V�h�����;��'        ���s"p8s)%����       `^r�B����ݑL`�<��1q���       p�D����TJ)V����'	�       8g)%�;0iw�3����K?gG�;       �̤�"�T{Ƭ�D�m�֞��G�3�s���ab��3        �I���R����;09�G�3�s��r)n�E����        8��Ƚ��S ^) ΄���p8Ԟ        �/p��׽D�Ţ�������ib�Zy����        ��}WWW�Z�j� ��]�4�X,�Hw       �y�Y�V�U����3��`�ڶ��r)n#w        .�r������3�&p����b�XԞq6��c��X{        �ȑȷ��}����w
T!p���R�}}�מrV��}�	        �1���.nnn"g�)pZ�u ff�XD�u�g��;       ��	��^۶q{{���S�"p���R�V�h�����$p       �7���G)%>|�m�֞\�� 3�s��z흐�H�       0�����R���D���� @�0q��X�V^|�����0Ԟ       �o�׼��R\__�j��=8sw�	k�F�~��       ����[�Vs�q    IDATquuU{p�� �u],���3.��       �<�Oc�X�������L�r����kϸw       ��,�Tڶ�>D)����x&���s���h�����1���       �L��\?�RJ|��!���=8#w��(��r��.�;1C�        0K)������rY{
p&T� ж�����nW{        oH�S�z������3�3�Y����c�X��H��       ΋����b���� ��3@%)�X�V�u]�)M�       p^���m����C�m[{
0Sw�
rαZ���R{�E;1C�        �1�{]9總���rY{
0Cw�k�6���3��       �'m�4��븾����x8��b�Ţ����       �<	ܧ�������RJ�)�Lx8��s�V�h۶���8���nk�        ���4M|��!���=��;�;k�&��w N��p�aj�        ���\q���R����z��=�8�� ���X.��g���       �7��4-����Ⴣ��7y�x9�X�V~�΄	�       �[J����i�����W_%pxcM��z���	�!v�]�        �#�������&��u�)�����b���rY{�!n       ��TN�r������Y�
��g�7�s��jm�֞��l6�'        p��yh�6�������`�� �m�X,�g���q��v[{        '�R�=��R�����.b�ړ�J� �(���"��S�������        N$�����i�xxx��~_{P����J)�^���3��ljO        ��r�J�M)%nooc�Z՞T���I}�G�u�g����m�	        �PJ)RJ1�c�)���jm�ƧO�\��mI ?(���J�>c��>�C�        ��K��<�m��G,��S�q��t]}�מ�o�l6�'        P��}�RJquu]���Ãk�p�\p�/W���������        *(�Ԟ��.>|�]�՞�#�;�7�m��ڋ�3����x<֞       @%�����s���������p��� �&�}�G�x�<'�ͦ�        *�9;�xF����m���!v�]�9�r��3/W���������        **�Ԟ����{ΒX8
N���׾ｈ=S��.�a�=       ��RJ1�c����k���nk�~��� ��X�V��3�z;        M�.��9���u��ܸ�3�O0p�rαZ�����Sxg�ͦ�        & �)��3xG]����Ţ��	܁������b���0�g        0�{���R\]]���Ffȳ4pQ����z]�y'�xzz�=       �	�_��m�?���z��ij 8��R,�hO{��x<�n��=       �	I)EJ)�q�=�Y.��u]<<<�~��=�oC�^�u�^�������7"        �C)��N�����q}}�?L��8[��X,^�\�����        ���R�	T��}t]�����lj��B����R�}m�֞BE��6�C�        LPJ)r�1C�)T�R����X,�������$�3w�t]]�y�%���T{        &p�i������v���>`"��Yh�&����s�)L�0~|        �*�)�Ǳ�*��>������x~~�=.�����R�}m�֞<>>֞        ���x<֞���b�^�b���������'�����R��m����S� �       �G�RbW�yUJ�����n�����P�����ib�XDJ��&ȋJ        ~FJI��?�}}����s<==����QJ��R{
���T{        3�r��f�\�b�����x~~�=.�����st]m�֞���������g        0#)��9�����R���X,����ݮ�$8kw`�RJ�u]t]W{
3���X{        3$p�G�R���&v�]<==��p�=	Β����R�m]�EJ��f�x<�f��=       ��9GJ)�q�=�x9ܺ�n���)��c�IpV���4M��B��O{||�        ����"7?�����>6�M<==�) �F��$4M}�Gι�fh�xzz�=       �sŝ_�X,�����#p�*�D��QJ�=�s�       ���s���X{3�R��r}����Sl6�ړ`��@���.����gG��       x��;�%�WWW�Z��������I圣�{a;o���)�a�=       �3!r�-�����2��������I�y/����'        pFr�1C��X{
g����?==�v��=	&Oi
���st]m�֞�zzz�nY        �TJ)rκ�T)%���_C��nW{L��x/a{�4�R�=�3���P{        g�w�K�4qss��!���]t���o�����{z||�.Y        ޅ+�i���:V�U<??�f��=	&C�
�	a;����X{        g�wN��WWW�\.c���f��9��S��E�N��       ��\q�J)�^�c�\���Sl�[�;K�
���i��(�Ԟ�1j�        ���Ω����*V�Ul6�x~~�����?�m��.rε�p�c��3        � ��SK�9V�U,����]7ť�ߕRz�SJ��p��q�����3        � �Wܩ&���2��el��x~~���P{�+�;�M9��.���3	�>}�.D        N�w������>v�]<??�~��=	ޅ���R�k�Sq<]o       �
Wܙ����8��lb����䬨W�WM�D�uQJ�=��ӧO�'        p���q1�Ii�&���b�Z�v��������,�mw�p)�h�6����R�9�U��!���k�        ����"�, frrα\.c�\���á�,�ew�P��h�6ڶ�=������        �R���I��>����~��&��m�I���pa����뢔R{
�/�        �
Wܙ����������[�B� ����*�T{���       ���ib���8����w�c�\�r���n��ϱ��kς%p�3�4M�mM�:�������        ��������.�������&6��7j0I�W83)��.����s�9�ˆa�����3        �J)1�8�Y*��z���j��.6����L����˵�RJ��jρ�v�         &���á��e)���>�����nc��Ӹpw���s�mmۊ�9+��.���k�        �o�9G�Y�Yx��^�c���v���nW{J�3�R�۵v87�8���}�        �]��;g�����66���sNJ�3QJy������)��}�        �])�(���x�=�\)%V�U�V��������q�=�3'p�	�9G�4�u]��jρww<�ӧO�g        �{��.�圽�]�ױ��b���n��=�3%p��I)�~!�9מ'�����}        f���á�xw)���>���ab���f��SxSw���SӶm4�?�\��f���        �i9�(��|�(9�X.��\.�x<�v���v���MI��D�M�D۶��@U�0����3        ���Rb�Ǳ�8�RJ�V�X�Vq8^c�ajOc��pB)��9�^jO)՞����'/d        ��RJ��3���i�i�X�ױ��_cwo��G	��}��R"�\{L�n������3        ��#���#���m�m۸����~���ew�K�� ����w!��_7�c���՞        o�i���v�g����/����|���HJ)��y�E��}���q<k�        �7�4M��3`���ݷ�m�v;�;!p������~�n������3        ���#�,օ��GD����ݛD.�"~R��o�ځ�7�c���՞        �i���v�g���Rb�Z�j������.v�]�����8!u.�����m�H)՞�w���        xWMӸB�����2��e�����v�Ǳ�<ޑ��"����x;��6���j�        �w�s��s�P{
�ZJ)�����#"�p8����Dr~��}�K)��9�ړ�,����j�        ��i�&�����������ib�Z�0���]w?#w.V���J{)%RJ�'�ٻ�����X{        ��K�����߮�������u���s1RJQJy��]i��z||��v[{        ��K��8$���m�mۈ��1���}f�-A;L��p�O�>՞        ՔRb�����)�����1����/�I���H)E��5j/�DJ��, "���b��3        ���ib��՞�/],!x�*�;��r���J;0=������k�        �Ih�&�C�@ާJ�l���v���R{���6k�        ���9G�Y8����p8�~����Xy�e�3I)���/Wځ�8�qwwW{        LN�4���c��S���A�q_c���ݟ�'pg����j�~�Ǐ��        ��%r�#�m�F۶�����8����;U|�������ދo        �)�h�&�C�)�oh�&�����+�/����c�?I�λJ)���8_��&k�        ��{9+~���+��0�����x���_�yS.��e;qwwW{        �F�4���c��S�w�s����������K����_�eĞs��R�Y@E�8��ݝ�        �^"w�r|�������x|��uyw��K��e�𥻻;/�       ��������BV��|-z����o���ߟ����H)�^`�<b�?���!6�M�        0[/��x�=��������%v���0�������{J�5dO)՞��v������3        `�J)1����T�4J)QJ��������/W��p�]�~f>��?�ʞR�o�p8�Ǐg�        �i����������i�h���/������?��<X�<Z��pJ�0��       ��D� o�{��0������͠�}�������� S1�c�����p�=        �NJ)ڶ�'�rt��m�~������������k����p��O�>�v��=        ��˕eG(�)�9G������c��/ÿ�����9��RJ1��߮���/}����\����x||�=        �^�9J)q<kO�)?¿x	��q�E���}��}D|5(�2<����q�j����n�q_{        \�R��c�s�y?������'>��p8�Ǐ��@        ���4M�;p~��; kq;        T�4��i�&� ��q㯿����P{
        \��mkO xww ��Ǐc��מ        /��;p�� |���]l���3        ���s�gM��W}��)���k�         � rΙ��xzz�����3        �o�9G)���7'p�o6�M���מ        |G)%r���ų �v�]����8���         ?�i�;pV<���>���/q;        ̌K��9�l@q;        �TJ)����R�) �M�p��c���1C�)        �oh�V�̞�����       ༈܁��\�����W���S        �7�4M�	 �L�p��a��?��p�=        xc)%�܁��\�a⯿���~_{
        �NRJ.��$p� �v        �/���D�p!�a�?��S�        D�̍�����á�        ��D�������x�       ��K)E�u�g |�����?~�        Ѷm��j� �&�;��:��?��?���kO        &"�$r&M�p��C���q<kO        &�i��YF
LOS{  o�%n���        `�RJQJ�����7 gd�ߋ�       ��R��i"�T{
�+�;����v�v        ৵m9KJ�i�lp6�M���_1�c�)        �5M#r&�3��=??��ݝ�        �-M�D)����5� ���ӧO�g         g��)�8�� �w������        o.�M�DJ�����03�8���]l6��S        �3�s��R����S��;�������        xw)�h��%w�� 3q8��?���nW{
        p!RJ�4��8�;�������?�p8Ԟ        \��K�9�N���� ���l6qww�8֞        \��i�x<��x�=8cw�	{||�����3         ""��!rލ�`��q����xzz�=        �oJ)�R���P{
p�� 3C|��1v�]�)         _�s��m�p8�8��� g$� ��9����       ��K)E۶�R�=8#.�L�v���?z7#        0+/�܇a�=8w�	x||�����3         ~I�41C��S����?{���F��atG&�1� z�C;օ�̌�~�&�r�\.I�I�$$߀��������OOOq<מ        ��p���{_{p�� +������X        �F)%6����mw�L�_�~�        pwJ)�K�� 7F���v�]����=        �Cm6�h�E��1P��	�>Ik-����x<�=        �S���X�E���;�'��9�~��ֵ�         |�RJl6�;�K� �p8����        ��UJ��v�V�B���|��Z�����pX{
        @
�8F)%�eY{
����,�OOO1���S         R�!��m,����� �����p���g?x        ��RJl�ۨ�F�u�9@"w�w�Z����8kO        �	�8�01���S�$� �`������W        �C�����K,����� +��K��>^^^֞        p�6�M��bY��� +���Zk<==��tZ{
        �]�!��m,����� +���������        ���R.��F���h����K���         ܵ�f��X�e�)�'�����OOOQk]{
        �C�!�|��<G�}�9�'����{�v���vkO        xH��6ZkQk�Ý���<�����-n         V6C�˲Dkm�9�����n���k�         ��f��֚åp�� �q�         �ab��F��5w�3w���{��n��n�)         ��R��{�5z�kOށ� "N�S<??��        pc�a�R�k�p'��C;_m���^�        p����;t
�M�<���OOOQk]{
         �`����K�Z�ap����i����k����=        �0�c�R������ ���x(��!^^^����         >�01C�Z��&t�!p²,�����i�)         |�qc�X�E�7@�ܵ�{�v���vkO        `%���n��Z�eY֞����[�4���s�Zמ        @�0ė/_bY�h��=��;pwj������q�)         $��l���V�;$#p�F�=v�]�p��m    IDAT��软=        ��J)��l��˲�=�w�.L����Qk]{
         7d��n���Cw�-�///1M��S         �Q�k��X�%z�kO��%pnRk-v�]�����         p'J)��n���V�;�@�ܜ���x}}�V0         |�ab���F�u�9�P��͘�)^__c�絧         � �q��������///q:�֞        ��)��f���{,����'�]�i�Z���5���S         xp���n��Z�Z��>��H����>���          He��!Zk�,��s��܁4z���c��	�        Hm��n��{w�ޑ�H�p8���K��֞         ���ryZkQk]{�<�;�������۴         p�J)1�c��V�^�_����)^__c�絧         ��(��f�G��,��~���T��)^__�t:�=         >�f���{�ֺ֢��w�S�        x4���1�a�Z��������        ��J)���Bw�9�;�!N�S�v���i�)         ��u��Z�Z�ړ �;�\l        ��+��8�1���#p��4M����<�=         n�9t�1�e���ړ`uw�_9����˲�=         n�f�G�[kuѝ�&p~��p��n'l        �wt��^k��Z��מ�J�����%l�6(         �qΡ{k-j�Bw���[��������}�        �O4C�R��.t�!܁�4�s���8kO        ��UJ�RJ�p	�[kkς!p�d�����1M��S         �+���l6Bw������Z������,��s         ��8��q	�{�+��O�nY�8���}c        �4�c���h����M�Ã:�N����x<�=         ��J)QJ�����;~����i���x������y�9         �(��f�G&\k�֚Н�!p�0�s�����p�
         �8�1�c��.d&p�;v��>M��S         ���0D���;�KFw�3�<��p����UV         �7J)�\u��
�IE�w���4��         ��ﯺ�Zמw�e�<���[�G��        ����U��k�Íi���p����X�e�9         ����{k-z�k����FL�t��         𑮯��ޣ��;�B������!��o
         �*J)����__uwٝ� p�dj���}Y���          \��0DD\���yOwH���4��p�i�֞         ��q�q#B�����Jz�q<E�         ��;���h�E�u�I�(�;|���7�ڽJ	         �'��;���>X�=N�S��8��Z[{         ���>v��F�݁`~J��:j?�         �����؝���;�_��i�֞         ��u��Z��!p����4��x�         �C�0DD�8��{���%z�1	���������         ��PJ�qcǈ�K��Z[y�I�����)��c�G_$         >�0����֕W����˲��t�i��t:��         Vt��q���%x??��;����/�/˲�$          ~���8FD\�����&p�a���͕v_�          nK)%J)��ױ{km�u��;���<�4M1MS�Zמ         �;������!��;w��~��>MS,˲�$          >����9zo�]r�s7Zk1�s�N��          g�0\����7��]x�A��ͺڧi�y�מ         ��(�D)��G��»�}=wnƲ,��}�gA;          ����{������;)��cY�8�N�,KL��ֵg         �@���s��{�&|�}	�I����e�y���         �4J)�����9t��������z�1�s�N�˅v��         �5���1""�q�ӕ�޻����Zk1�s,�r��.f         ����{D|���N�λ9�����          �u�.�������˲\.����<��
          ~�_]z���{km�����S�<G�����          ��r��Ϯ��?B�.p'Zk�����GW�         `=��ޯ�c��ϯ}����~	׿����          p�~t�����־����H��O��ϲ,k�          >�9|��~��3^~�߈���=           g�������:|�G)��#x�{��h������[yK           �v�R.��G�������s�~~j��{���	�         �[�w��u��� ��bx��w���Zkߜ�?����w�#v          �Gv��j_J��O��?�G�����~T���������Z��          ��q��o!p�߷���g           ����           @��          �$�           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���     �?v�ض�0����Q�EI�:l��>��H�3b	����@(�lŏR���7���     $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p          ��\�    IDAT A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	���Y��ײ,��; x����g  \��t<��\fY�׻����  ������t:����̲,���� p-��Y���P��_������l�� ��0�����?��\��������  ײ������m��2�����u�2{ ��l��7777��w ���           ���          ��          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�      ��޽=�}�w��>���@K�C�q:@ð	��a�
�)�7�E۸jS؁i;�%z�ZnI�~U���W�VK�np�R��.T\�2Tͅ&$)3$!�p�p>��i-�g_D�(	ؖ����ݯ�_�QI��|   @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��; {JJ��Kw  l��rΟ*\�����P� `�|��j}�tp�r��,� �r��}zzz\���&� �����^�j�n��w真]� �}'�|�h4���ѣ?(l��s���oI)����� �&���8���q��k��%��ׯ�o�9/D�o�� �D��8�R�Å��A���=k0��ٳgoJ)����� x�����'�c�+��뽱��["����=  O`�s�'���C�c�+���9"F��#�U8 ��<�R�w4�>|�k�c �t� �y�����ht]ι�Z� �"9">�st:�SJ�t�}z�ދSJ7��n���� ��0"NE�j���|�`{?~�U9���K� @�|%�>55�>??�H� �>w �ȅ��,Fā��$ P�و�����v��w�c������mnn���J�  {ڷs��Vk�n�X:(�رc�LMM�+"���9 ���pJi���q���q� .�� ����oH)�AD�3"�Y� �3��R��x<,..~�t�,u]W���RJ#⭥{ �=�3���p����R:h��������sΝ�x}� `ϘD���dr���o?S:��e� O�ĉ/�F�\��B� `��bD�UUuw���,4���ʛr��q}D\U� ؕ&�ɜ����Y�`g�R. �6"⾔�����J� pe�� ���`p�h4�n2�N)��t �;���L&��N��`J)��v���՗���_u^� `W8�GıN���1�����^�j�n�9�'"�U� ���s�{<�<r�ȏJ� pe��%�뺚�����ҡ����= ��t.">ZU�r�����1���oss�X���X� ؑ��s�+�tg���~�`wX^^~aD�x�(���{ ��'���8�o߾����F�{ �� �4�z�7VUՎ��#��= @��8���R��n�t�;]8�=PU�b����� v����������no��v�����s�="^W� h�ID��9��v���`���e��z/N)ݜR�-"�_� h�/Eĝ��𞺮/��~�ڈ8��9 @ä��L&��N��`J)�����s���o��RY  ��aD����N����1 ��E �"kkk�677o��vD��t PVJ�LD����y`vv�|�`�Z^^~eUUs9繈xn� ���qι��v?[:��VVV~-����Έxf� ��o��G��G��A� �3p�-V�u5==} �t0"�Z� �V���X�y����E���---�o�Z7E�|D��t �}r�߫����x������= ;q�ċF��-)�[#��{ �m���x�p8�H]�?)@s�����~����F�;"b�t p�<�R�7"��\:��\t�{$"~�t pE}1"ֆ��=u]?^:����G��u���pJ鵥{ �+&G�'r΃N��`J)��y�`����d<�]����J�  [�#b�s�@��}�t������Fġ��!"Z�s �-�R:3�L��E���K� �k����#�X���\� ��� ������V�uSD�G��K�  O��)����̟��Ξ/p�VWWy2��9�^DL�� ��s��X�t:U:`+����)�<�G�U�{ ���9������t:�/��`� \�����ۥ{ ��d�s���v��t��0�s�ܹ#b!"fJ�  OɏSJ��ˋ��_/p%�z���nN)��/� <%_���UUuw���,��b� ����k#�PD�#"�
�  ��FJ�C9��N童c �����U���m9煈���= ���券#���n��X�����oss�hG�kJ�  �^J��d2Y�t:��r� v&w h����WVU5�s�9"�)� �?��Z����t@)�~��q0"���9 �祔�D�ə��fggϗ�(ᢗrF�[K�  q.">�s�u��ϖ�`�3p���9w�܍)�v���J� ��pJi���q���q���8~���rηEĻs��.� {�(">�R:�����1 M�\ ('�����>�R���n�t ���; 4����U���m9�vD�f� ��&q:�|���>T:�Ɏ;v���Ի"�/+� �ݣ)�{G����Ç�V:��VWW_1�Ln�9�E�sK� �.����s8�S���c �}�`���o������h���d�Ο?|qq�J� �$u]?c�����;���= ��|%�>55�>??�H���diii�պ)"�#��{ `7I)����333��Ξ/���e� ;H����V�u0��{1]� v�o��[�֠�n��t�Nw�(w1"��s���pJi���q���q������jzz�@J�HD�V� ���E�ǫ����,����M �;v용��wED'"�C� �I�gJ�ľ}�����mz�ޫ[�֭9��DĳJ� �1���)�?^XX��c v�~�mD���K� �T�8����x�������1 �-� ���u�����_�s^��7�����D����n��P���`yy��qcJ�`D��t 4�FJ�C9��N童c �����_�L&��� O��qG���n���1 �M� �K���7G�bD�@D�و���j�����ߗ�؋��գ�躜����= ���9�=�O9r�G�c ���`�s���1S� � �t&"N���<0;;{�t {�� �2�^�խV�ֈxw��٥{ ������Fw=z��c ��r��RJ�������� b}}���p��/��F� (`�SJ�����1 �S~� ��`0�ųg�ޔR:/-� ��#�}���#u]��t ?����RJg���+l�s�'���C�c ��.����GD�p \i�����F+��Z� ���`�W�F��r�݈���= ��rD|"�<�t:��r�  ��'N�h4�ra���{ `�#�TD�v:�ϗ��;~���rη��r؝��s^���Z����t �<� ��\���bD� `g;�WU��n���t O�EG����������z���������;v��5SSSnD��p \��SJ����Su]�K� ��1l�=hyy����Έxf� ��M)}h<�Y:��S�u5==�;)�C�{ �}&���o߾����F�c �:u]?c�����;���= p	&qz2�����ϔ��Ka� {؉'^4�n�0v���= ��kUU��n�7K� pe�z�7VUuK8���&�ɜ����Y� �</��ClD�})�����/�����\ @��G��u���pJ鵥{ �RJg&��R��y0��K� ��z�ދSJ7��n������F��q���|�t ۯ�뽺�jݚs~OD<�t \�������#G~T: .��; ��u]MOO�NJ�PD�n� ��s�Ѫ�����ߖ������}���7D�|D���= �Y��9ߕR����|�t �-//�0"nL)�����`oJ)}:"N�۷ﾹ��Q� �
� ������XUU;"����J� �'�8���R��n�t �s�(�����[K� �g�MD�UU�'�v{�t ��ӗrsηG��J� �'L"�t��d��}�t l5w �	�z���nN)��/�������s8�S���c �z�ޯWU�ވxGDL��`�I)��L&K�N���R.�@��S��˅�r�M [o�"b���|�t \)~� �����}���7DD;"^S���/�t&"N���<0;;{�t ;����K���܅��?�t ;�و�?���v��-�ε���k9�ߏ�wF�3K� ��};�>��8z��J� ��f� \��������#o-���3����W���_��`�XZZ��j�n���F�+
� ��䜿WU����c�T8    IDAT`qq�{ �=N�8��htKJ�ֈxA� v��D�����G��I� �.� �����~����F�;"b�t ��hJ�ވ�/,,�s� v���VU��s���{ h�/F��p8�����K� �{��G��u���pJ鵥{ h���9:�΃)�\: ���; p�VWW_2��.|��y�{ h���A���n���1 �-�~�ڈ8�r�7RJg&�ɒ� ��K� <��qD�t:�+ %� [fiii�պ)"�#��{ (���`ff�Ogggϗ�`o[^^~eUUs9繈xn� �9���N��W�c `ee�M9����>"�*�@1��9�?�tg���~� hw `�]�����ۥ{ �6��8�s��n���c ���9w�܍)�v���J� �m~�R��x<^^\\�z� ��z�ދSJ7��n����`�|!"�WU���v{�t 4��; pE���k#�PD�#"�
� pel��>�s>��t�Z: ��EG�G#�7K� p�|9"��9���>V: ����ھ���"��)����R:3�L�:�΃)�\� ��� ���˯��j.�|sD\S��-�O9绦������) OG��sD���GD�p [ �t&"N���<0;;{�t \���rF�[K� �%�E�Gsνn����1 �t� ���9w�܍)�v���J� �<�Rlll���z\: �B����V�u0��{1]��K6������/,,|�t l/��l9��UU�����v��{ `�0p �X__�j8�-�܎��,����D����n��P� �R�;v���Ի"b!"f
� ��M)�;�V>���1 p�����b2�ܜs������I})"����u�x� �i�������#�`D�="Z�s �׆q�������t l��������+�܉��R���+9���������GJ� �vYZZ��j�n����xy� ���ҙ�8933�������= �S� ����~��j�9�^DL���㾝s^o�Z�v����1 P��\�Fy8�4���8U���t �R�u5==} �t$"~�t�w.">^UU��n�e� ����9v��5SSSND���9 {��L)�طo�}sss��1 �$ǏU����xw��٥{ ��ID�N)������( M������CqC8��N?N)}x<//..~�t �&� @c�u�����_�s^��7����&�ɜ����Y� h��`��gϞ�)�t[D��t�.��R�P��x���j� h����_�L&���p�}9"��9���>V: v#w `G���o��ň8��U�F���V������t �4�v"���{ v�o����'�9��1 ����;w�ƈX����= �EJ�LD����y`vv�|� �͌� ���뽺�j���9?�t�����]��莣G���t ��r._J��qrcc�T]���= �ӭ��_5�v���(��CM"�tJ�>U: �
�h v��`��gϞ�)�t0"^Z�`���x�p8�H]�?) �������?�9�'"�U�`�D����n��P� ح.����GD�p�N�hJ���h�r��ᯕ����� ����գ�躜s7"~�t@��D�y��tL)��A �,//�0"nL)�����h�aD����N����1 �W?~�U9���K� ?�Wr��SSS���󏔎���� �5.|}d1"�� ������Zj��W: ����ro��ו�h�o��[�֠�n��t �Uǎ�fjj�]э���h��SJ����Su]�K� �^g� �:���oH)�AD����= ��)��������7K�  �"����[.|��Q.�}&���o߾����F�c �Q��3���}ι�/���&qz2�����ϔ� �7�D v�'N�h4�ra���{ ��/F�ZUUw�����1 �Ϸ���k9�ߏ�wF�3K� \A���d�y��v��t �ļ��!q_Jieaa��c ��$ ��7��F�M&��)�ז��J)�3��d���<�Rʥ{ ���[#��{ ��و�?"�u:�ϕ� .M��{u�պ5����R.��|+�|�x<>y�ȑ�� ~>w `Ϩ뺚�����ҡ����= ��\D|����v����c ���(�E��s�+�tg���~� ��,//�0"nL)�����x�RJ�������onnnT� xr� ������XUU;"����J� <E?N)}8��k���( l-G���7�VU՟�����1 ����Qn����x]���h�s�'���C�c �Kc� �i�^��)��SJ�E��K� �_��;���=u]?^: ��VVVޔs�G�@����L&��N��`J)�� ���s���o�p�{ lN�fFĩ�X�t:�/ <=~�  �����}���7DD;"^S� �_�"qrff�����{ ���(h��qι��v?[: (cee��rοg����o��G��G��A� ��� \���jzz�@J�`D��t�'�"�c9�n���c �fp���s�^UU�ǃ���o�� ��ĉ/�F���n�������D�����G��I� `k� ��^�׫�zoD�#"�J� �ޣ)�{#�����ϥc �fr��ňX���u�x� ����գ���dr8����=���#�9�A��y0��K [�� �I����d<�]�<�t���cDr��v���� v�~�mD
G���R:3�L��E �K�(���F��q���|�t p�� <EKKK�[��M1//��x��333:;;{�t �s����b2�ܜs�o�(�<�"�����t��t ������)�<�G�U�{��9������t:�/ \y�  �袯����.��(��8�s��n���c ���Q.p~�R��x<^^\\�z� `w��z/N)ݜR�-"�_��Q�﫪��v��Y: �>�  ����_�"�1U8h���҇r��;��WK�  ���\�|9"��9���>V: ������mnn��xM���RJg&��R��y0��K�  ��� `,//��������qM��1�)�|��������#�c ���Q.𳤔�D�ə��fggϗ� ����rF�[K� �q.">�s�u��ϖ� �2p �B���9�Ν�1���9�R����SJ����Su]�K�  \t�;�-�1������/,,|�t @��\ "�����>�R���n�t ��  W����U���m9�vD�f�`[L"�t��d��}�t ���(��GSJ��F��Ç�t �ϲ�����dr��\�S�w��{�~�t �,�  WX��sD���GD�p���q�������t �S�(����ק������) �T,--�o�Z7E�|D��t��RJg"���������K�  �d� �Mz�ޯ�Z��9�[#�*�\�����V�5h��?, �t]8��F��Y���K)-mll���z\: ��뺚��>�R:�\��<)��s�������,� 4��; �6�����tpyRJ������[� `+,//�0�������9����~�t �VX^^~OJ������9���z� x�|9 `�yjv���?�      O"��u) ���          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��           4��;           �`�          @#�          ��     ����An�0 AP������0��s	��6S������Y     ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           �88C  �IDAT$�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $� �s��g       X��� ��E� ��qow�       ����  ߋ� `�9珻g       X�w ��; �zw����X     ��s�S .� ��/�`�y��{    ��Y4�p?
 \"p Xl��l`��{    ���9��x
� p�� �b����w    �������Ш �8<  �g�;l�w    ��u����Q .qx  X�w؃�  �c��{ �g9�S�ch� �K  �s��1~�=  �ߎ�x�{ �g���a�9� �^�U  �9��<� �6��|�{�9朞g `'�60�� �2  �� �0�t� l��xba����g `���܏ W	� �� �0��{
 �������3 ����"p �1�� �H� ���6p��h �Ɯ��61���
 ��;l�0 �?�SkJ+�?�    IEND�B`�PK
     ��/Zp&ر  �  /   images/aaaf988e-4d8d-46a5-ae55-a0506af48a51.png�PNG

   IHDR   d   �   �K�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  >IDATx��]{�T��f��{�e��"b4V\QJTb��jbI�ӴZ�4��F�4*R�IM�Ҵ�hl�?L6���
ۚ(�y������;;����W�߹�w����̝�z~ɗ��8���~����{*��;wҎ;hɒ%�D(�N��H�R��� ��x<N�p�B����bŊ�$d ===���d2�}��qR �E���d�YgĹ�~)y	�d ����F���k���Ou�r!\�/M$7�����͛����ܗ�;�E�
�̟�ȗE3R��dl��o�$�!`!2�X^�>5�a9��,w��q����ŤQ�����($)����X�#�jb��� %C��:ֳ|�4j�gY�Y��A���{X$Oa5�s]
�������b�U�U��(��v�do�ǐ�Y���n�q��� �~He0C��s�|��%!��P��.$���Ç�F���Iss3q�=��I��n�U�188H��:*�V4��ҧ$��yb0���W�i2�C2�̐�$$+ڀ$طoMOO�3/�2�ʝH$��������n��ۻw/MNNj2��g跡�!s�p���~��T�FY&X�XRd�&T�V�Y,��(�� ��a!�䊒�)˻,��e9�&���P�@Eќ\�r�R���b�������S����h�*F�z0��W�]d*�`-#,�Y�k�@ЗYnc��h�����)a)�tV��;t�J1�#�M,��u��իf�q�F�B�a�Lr ��ycvh6��6v��Ms��U��7��s�_�L�/�=���3������7l�`?<��S�gX�`��C/�����,x��I�����,�-d>O=����a�!��Y�#�c��xP�ӇO��'�"4�7���U�����Y��ʰ��u#�k�)*���G��8�@��L}��-��}�M�I2�H��2$�`4u˖Z?�߄�usD�E���n.���{,7��|#�[u	����u�H\�t)����Qt����7�r��7B�����aBĂ��{L�߀��tv�9��͓�芉�I1�Z���o��*�G���f�V��7�m�|�NM�c�iin����3�ې�,ג�s��;�[���SSccM��B>y>��d�ÉZ���k�9k��ɶأ������/ay��;d��f�&1� n's�mfJ��K�|sY9H���M2\<#OV��D`]�/X~케	�Z�7B0̏ye1��x���,���[�� ]9M�$���\2����΋���j	�����z����L&Apg���1ഖ\֓� ���YV�\��T�䁐@�|#���o�d	��AΫ,�9m�Q=�����9'�$�f������
 �g"�
����׋Y2�M��Y>d���1�Ӵ (�6�ա=̧c`�\2We.�>;�2��:O���Ԅ���B0�/W^��<K��0W�xR������&���E��.&G�/�3���0�+?��N�Ƚa�������)������}&į�Je`I�$�ր�Ѹ�;~�|�v(A�,���Z,��j��3����ePJ��{�G)��j#��E҉�!Jr9A֤)G ׺��"�)w����}�g|bBLBG"�~FP��7j"E������Hr$�k+���Z��R,��([\���(Mr�GZ^0��Zl�	�C��(_�"?!��@``@g�F<�^�r�4��8m�
u�S��C�����S��a��p�I�i{�?�qZZșM�bЄ(M�bЄ(M�b0N�f��$�ԛ�-BR�=�+�5�SP��+��B�����j�n�:sPP�:�(��R�Š	Q�Š	Q�Š	Q�Š	Q�Š	QFP��W)G����(|�100`?�C�>C�Š	Q�Š	Q�Š	Q�Š	Q�Š	Q��E=��3���.�k!����Bl�h�C�tPW�ⴵ@��K�;r�W��������)!F ���@I��!���ܙ���%�M'�����P�8%�t��B�@͡$-�? �K���9��.���愩!�����94�T�]:;Bu�T��h��m��h�x�Ѭ1:�y���Hsd��z��2��i��%m#�����iW��K��BP7[�#hJ��#���|�HKPS(%��H\��Fη�Hf��lW2B�Y=��Y��3!Υ(�B��`��-�u��,7)(�>�ݫb<tY��h3���q.eS�[�ӧ��Rv�̦���4����#4�1F��F�l��R�N6��$y���Z��dKN7�|�Sf'�l���g���q��S�����q_�&�∧1$E��g��U�� ϙ���s�g���X�y"�D�̽1�5��r>��Mp:'!�4(�:��V�d+6�'�ژ���=gO�CNq���ɹ��n��ΰ0���(��~ܻ�N�r�A�r~`�N����X�+�n炖qZД�r}(�S��ge��9����t5Nѥl��������#�Պ!x��x%B���muٯ|������u"��i��I�)R��2��d�
���������`������e�;���-6��eA9v?�r(&��R�<s-]����0_����>c�X�$��x���pl	��bc\9�=���5���.���5b���/=B�z���*x������r�V7�V���P�#�^�,+1Y�~��ψ3p����j�SB��G���X��n��0HS9���J��;���U}0�ε������m��:f$ZF��чl)}l	�j���L���ܻ1��c��VfK0[[c��q�3��y,+��A�sI�ZTOM��p-B��7ZF�p�=7h�k���X�95�$��q��ץ{s.��y���:s�{lqF6�s=[���˂�a�osO<�	�q�T2����!k%��YY8F���D+����&��9f�q��̀6�MY�e�������Pz����Z̅��X
j��r���XJ1��y}��{�"`�gH�;ŤOHY�JP���r	p���(���b�4}9��!�A�4!�A�W�(m!�A�4!�@�j���B8����MR4�I��7v§���̅���8k[!�J��b:� ���Wؔ �4Ნ
�d�`�4\C�&�2�����\�,C�;��M?6~<S��@F���*����ޤ�i���D\�]r+�hR��-@Y�^���n��
6;pKP!�2�h��U�cF)(��D���������RP!2�ONN
ץ_����466�����iSQ�4��U�ZP��7�I�����A:����^;ؖ{��m�5��^Y[[[����ݼ�ط�F3VaL�����_ �'	hjj����B�E��T��Dn�V�h����0��(�P*:�na- ��ikkq��a����i�.�;H����� �R�ݻ$�"����s_r{"g�`txxX|j2�C��;c�]��+��s@{Z[Fy������˲�p*��T�*4�C�/�ru{�����fǱ�L��	@���t_��� ��ϩKh��.�~��2�1A�/�2 Š	Q�Š	Q�Š	Q�Š	Q�Š	Q���/�d�O�L-�	IH64,�,�D:
5ttt,$�0�L&����G�\�e�WiY֌��u$�=\V��ٳ�À+U�]�Be�|��Z��3������?��emmm;���*D:�~�������5�yf)���?�v�ڞ����|��=E�ڻiӦkFFFҝ��3��縐���=(�w˖-W�۷/����2�W��������#. ��2��-���&��|�Iօ{ｗ�:�,O�b�c�/���ެ�V����+�ӻw�._������*�����R�ϟ��+/��˖-.e���Y,X�uY�r�J1��}����.�*O�ڰa�xW�֭[]ݯ[Y�A�4!��B��=z�b��,����꽯%?s%�����,s�r|^d.k��,]�5P�`�*�ۋ����^f%�b���.��Y�)#�wX�a�
����e,w�������޵�z	* ��WY堼�e����Y�����lB������GX~�r�OX.+�L|��i�c�����������>ʲ��V���Eʚf�'�o��LY�ȷ��O�l��u����Ye��[��KY����~�z�8M��9��,o�\S 9F�ϰ+���p������Z�:���z���|y�(�E{�(���z�*�UY�P���Y�&���P+F�$=a?p��9�E5.k�H����'�^n{�b-��Ls����,	�Q�Š	Q�Š	Q�Š	Q�Š	Q��Tx���� ��    IEND�B`�PK
     ��/Z��[.�	  �	  /   images/e8fbe2d9-26e0-4ccf-9f9e-bb43371c63c2.png�PNG

   IHDR  !     ����   sRGB��,   gAMA  ���a   3PLTE   ;;;777333///111555999888---,,,000:::222666...444hhPF   tRNS @��f   	pHYs  �  ��+  	IDATx^��ao��E�!$JH��m��JG�:C�~Stt�����e�ߎ�8��8��8��8��8��8��8��8��8��8��8��8��8��8���w7p������K�,,]��_y��6�]})���K��	=��R*K�z��6�]})���K}�$�->}p��T�.u�3��gW_Jea�RO�U��珮����ҥ�~�A���՗RYX���O<��\{-���k=��}��&��/{B�>��Q/7y���'����6�Я{B���v}��S�W>�7��n�"�Jea黧���~�Ǉ7��n�-�;��%����������7|X��s�_T�� ��K?��}��=�;���o>~�����O�?vD/��z}�����?��+^�?�U���oBea�?|ż\��}z���������O��k�P������VB�,,}s�	�������Gw+*K߼�˿���?�=��3zy����ϩ,,}s���Ɨ�~�Ӈ/���q���Ç����'����S>_y�?=�>���Nz�x}���'��.�<>�~y���×��[?~�SYX�������۾��N*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*���U*K�T�V�,,�RYXZ����Jeai����*��q�q�q�q�q�q�q�q�q�q�q�q�ql���)�Z�`�K    IEND�B`�PK
     ��/Z��`  `  /   images/95d79837-2dff-4c75-b12d-e13dc3081ed5.png�PNG

   IHDR  !     ����   gAMA  ���a   PLTE   ,,,444;;;�lZ�   tRNS ����-@�   	pHYs  �  ��+  �IDATx���An!A[����f���Uu�G��              8bx?31E��PQ�\Z�a��%��'Э��%Y�PQ��Z�I��!
�k}�hh�B��B�&���P)�^[�^h�о�7�_h�h���>��ޭP:���Dk���*���К�~����9�X�����C}�����Gy����;��*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ�(T*
��BE��PQ��            ����'{��˻    IEND�B`�PK
     ��/Z�l: : /   images/bce349f0-9fdd-490b-ade4-f6d95f909232.png�PNG

   IHDR  q   �   ���d   sRGB ���    IDATx^�}x]ՙ�:�ޫbٲ�0`p�zoI^����MI�������!e2I&$B
�3nءf�'eH���S\�v�i�}���HW�`[�-�����k]�������_�o�l��A� `0#kĵ�4� `0��A �ę�� `0��D����i����A� `0�3πA� `0���!q#��L���A� `0g���A� `0#C�F`��&��A� `0$�<��A� `0F �č�N3M6��A� `H�y��A� `0�@���f�l0��A��8���A� `�7;�4� `0��!q�0��A� 00$nv�i�A� `0C��3`0��A`"`H��4�d��A� `0�ęg� `0��D����i����A� `0�3πA� `0���!q#��L���A� `0g���A� `0#C�F`��&��A� `0$�<��A� `0F �č�N3M6��A� `H�y�p����]��X��S*��z�m�P*M�B���-�J�R�eY���R
 ?�e����
X�l�?z?�?MS�ݲ �]�*��oz�m>����WS��웝G�Ԫ�Aڕ���d-�R���o�ݳ϶���}I;{������h�1#i�|�]W�g����4EXI}�Wvof;��f8�c�>x%�}�����Je��#W��W�e��}�{��>;r����3�3�������6��h�m�}����mm�<�Z���O;{����ϱ��<���q���{_=��>3���S������c�n���8�;n�oz�~����X6����l}^��j�l8�=F*�R�,�w��x���v�<Hr��߲{�,˵,�SJy�	=|%˲ڔR+�0|䢋.j���1��l����˭�F/^���}��o�<�@��
Q9�m�tq��ѭF�d�]4���ĶK�v���v����?w��'��M�v���v�]}Wz��`��=,rΑt�`�����`\����@����_m�_�������ڹ��#������=��ذ-�\�kǥR��R�,��~z�u�ݺ�1����w�@i/��+Vx�}��ʇ.���$��8��Q*���^|������E���$��M�:-Z���s�~e�ލi�@0$n ��E�,_�z�K�������jUZ�r��(�,q{��[1{i!�]�6��;�q�5���;���Ŏ"`H܎"���jժ#�k���>򑏜�8��!�-�i�3�A� `0/-GK��k�2��W_}�?�V���n�����\�r撻����_~,-qi#�ˈ�0��j��p}�'}�_ �J0hP�]}>���`� �e����Q)�&�p������A`/B�Ͽ�D�T����|o,y���e�߳͒���[�{W���M���eAg��|屵7��+V��=�]��8zL�n݊�o���k���3C�&s�=����a{��抃� Iܢ;���c��,$q��!��A���[�S��[��S�� ��T�9(ˑ{t��W�w �*��*����|��I���P����-��I�Z
~X�gY�Z���NH����%�ۜ�r'����E��*vR8I��(�e{��PU�$��"xV(�R��&�$������~��5�U�'%��}��U{�T�2�6Nd�רZϸQ�?��ذ-W��wW��\[BMT����� �������ڰp��ν��ҩ�iF�č���]�|���.Yz��?��X�T��.����v�rà�N�*�,a�I�cCb��WhhB%Ls �=}oiR7��d��i�D��N �S���=[��K]$���!�BՉa�

�"����� �T��Ɇ��# !q�K�������	]�OY��PV���{J$ov�%\�w��&s��	���I_�_k$M���SY�q�Ȟ�%\�ZH��c!�C�<	����qR��|�I܂�=o��O���7MD�D0G⩖/_>yɒ�n����.�\��K��$?�y��sKVД��\O<��=�4:��h�K_���ObӚK�����vy��$J��1�7q�I����<�MQ���I�c���f3�,(���ʆ� m���S/'@�j���i����CR#^�X�]!l
�<���@�Q��f���7�~�Ӕ-#tB�j�
#.� [���ea��V�1���8!}�
�%n(P^�4$nx��o���??������?��1ˉ8&6p�����H�Jc؎'�p9��h�]X�d)ֵmF.(����c6�k�Neir�[>�0����Sp�2�9�o���Q�V�=��>i������0��0$e���2���UU��t�XVNPQ�j��$��2�%��H|�\�$b���w��Na����o�7���<o�E\i��k�H.�q�'3�MÜ���FW{B7�0|r����7̛w������k7H�?��C������R��Z�څBA���/ѯ:�v��Oi���뿧0�H��>���?��R�D������qsss�y�椫�K�u�Y�����/�zv�3s/�s�E��e�p� ���ʳ=׳�Dq�EK���;�b�歰�TiA�k��C�B�ڴĥ� *$��VLvc�a	�-��Z���\����>�A=��>�6���}������-������]1�� 7����%�+�r�Y#�rd�J�شz����$�;�g!����~z_+� 	�ili�K�D�GϜ�_:G͘
$�!q����W�5��k_�g���W��ը%K�|�����0����0$;PͭK��_<mK�������Q��J@�\��(��?R��N(۶]UJu[�ծ�**���㍚0a�㮾���I�H�f	Z䆻�Ȏ��D�ea1I�ҥh��)��T�x��8���N%1b�|k��z@�+�0�"�U��X��F���Ƅr�+�rF�_�2'���vs�A`(���>��,qqgG�'"U�	�`���;$�
I-�[{S��
��LI��Q���l�!�l-u��H��S��r�B��9	��:�9u
�\�AL�rW��NH��ĸ��.\�m�ذ;���63� �ˢE��������D��$AtE���ʭ�T���
`K����N=m�W����K�Y�(9"���x���*�����n_��,�֮Re˽�2���^���h��FAZK��#�u��Y�D��<$�|N��T�3�6�� ��J����Y=��p'����0M��B�*i��+������
��ڈ�f�����5S�&�m��q�D�ń�^��+�#��b�C�����6��XVyw{�`�l����,��I m�iS����Qӧ³�����wx�C"�Qu$.]�`��&�a�X��#���[�x�o~󛋢(�ƗY��%�f�����"!��)��i��f_{�=i���b�H����-X^NH��_��bYdFXn~W6)i�)�.ۍ��ø8-1��hn�
A��	V�3�5� ��J{�Dҷ����w���k�ݛ`Ȇ�r��%��X�5�S���kD5ܚ�b����Vn-7BFJח�qa�e~�:�V#q��(L�$��4I�P�Θ=��q�"$/�98�C��K�`挩��v�J���E؞"r�$n���̝{է��'���+0$n���θ馛uuuY�	�N9�|�_ԺGu+ʑ׿��K��bY}�H,���/Ŧ��'�n����<�E�xVs�p��@|�
U�1�Ι0
B�+uhK�N�L�3}e�n��y�l��
y[R��D��b��\�hk7<Sj�Hl.�h������Y8�w�*F�2Y+��Eq� 'ކb�� W���auu��2o�[cq�Μ~.�33�Ma�����c箌);�K5����t���Λw�'v�x��G���A��ŋϼ��7`��)�G�,�w�98$.s����h�����$t�XQ�9 �K#��Vp�~M8�cly� I\=X�����d��Y'�;���y�,U�ŲB�#�s!q:k�/���_r?!q6�8E�Hk��r�|^�޴�1$DB&�fY�f���'N�t[����+��#�;j��|�L�6����K,X��y���.�����!q��a���?�[n�%n����8E򖝢�%��Z�-E[{��ĉ���_����ZN�&1::k�J3��qaZ�B���8{�(��@7PK�&z��� =�ip��K���x�V���HH\��#�!qdm�,��ZTgcb�+��a�,��%�+ww�W��!/	Z$k�������b��k����՗��]�1+���1fL?�Ϟ]#qڵ;Ԗ�M�6%,��ܹW~l ç9d#0��k��`7}��ųj����ltw�|�E����C��%�K�zs�(>�u���kI��H��I�V����K�Z��b�6K�մ�ǷC|��@���f�ێ=7C����Z�j��z,q���Q�@�g�$��,�W�x�̠��.A໠ͭ����d�4�(�-�w]�2�|�o�=b����%Y��c-鉖��N���_��y������f��C��'�ϟ�-��Bw�a���;q���e�d�� e��Yѧ?����)�z-�+�AG�'/e�ݩ�~�&qb��T�11�R�Y���c*b�S�.�Mk�ᲀ���Ԋ��q�S�gp�8dnL�I�<���;��B����8I\P���T��{��o슎T!��(��Y
���8j�tq�2��F���������U@�L�WW�Yg��f��ҝz�p�ĩ�p��+/߉��� �+��^p��s�-:��o\���}�!q��鎞eGH��Z���;����8+��4��@����{�GR���ZTԉ�ΔNl�Z)��4��5w*��$8���b�^�ɍm��I�]]	���A�gEZ���/߳�0��4I-%
^އga��Lׂ/^sfs��0�����?]5�X!���õk$�OR��v�\��s�@,�:���Zb��C�N��\�B[[�^K�}�і�˗�0�|߷Ǳ�$��ժ��S�>�c������o����ʿ�'MS�M_���|�7~ǿSL�u�Ĳ�
�N��^�袋j������5��b�[3���o��]]]��۳��=G�-q�$n��%���%.�jJ����zf���S�'�,;��\�9�pA>�E�g�6W3|wb�?$L9<ٸ�3�SU�l;R)a�ک.R�!,�E�_m)����a����)�����/�رMB��a"�]%\��/�Ǟ��jW�X�z��z�o�$.K1�i�ӏ��\,��C��ZG�`���ϝ{�G���<�OK�,9����׿���R�t�Ѿ��$oa�do��:$\,V��,�{���{�:R���}f�ՠ�H�2$��}��@Ѳ�N=��o}�k_��Pa�Z�5$nzŐ�A q���q��6K,q�B��Ɯ1֮&4�<!qR�ڝ�,:��WZ☝ZK����w%;�5���9� �G�%qR+����{:S<U�Pr�N���v�}ҵPi������$�ĶE�N4�\�x����#�?�,��]f>���UN���?���~Mo�k�j]9}�٧�ok����q�Zv�%c��)`��PZ��:	��8,Xp��s�]��=�y�|�+V������?��O����S�0< M�I�mO�˴Ki$a��<���	��_.�K��~��������WJ��쌆��>G�'q=�:k>�p��v�TY8��SE'.��3�vۅ�ę�g6�f��
,�8�S�N�歝b��2�z�SӅ��ǸZ砡��y<���Y��q\��M��eW��\T��x[$F���TUk#ڝJ�-w�(ě� �#�����1q�����]��ک%�'IB�z�c��� ����A��b��ɸ�s�ӎ<���@W)F����˞Y��b.6o�2|L6��S�u[7Z4���8y��W�N����cI�M�̝j#Q�h�mX���������n�̢E�Ol���v���a
��I����ܺbŲi˖-;cժU�b��y�8��$Y�@�b�b��Q;�����o|�g�}��4�5@0$n�C��]>ū�8�SI�B�o��2�m!�"	�f6�\h��v}l��	شƹ�|���/�R6�~�*�Р�S���F�BC�v���	F.�t�Nl�$Ε���k#q���Z�2XR���:�դ.I]�JUq���|.z��1���TC�������6�曾�����p� �8�'��������7k�j�T~�ڭ)�Ϙ�������*C#1B�#Ua6����񳅟���>dM��8.�z܌?l��Uߠ�ZpK5���ƶ���{�e�e��V��G�u��Ìj�s����~r����y'p[��:��{ZӜ\U[,˒�������4�eG߈W��:�D��N�����y���(�#l?C�C��ĉC�
�G�q
hi���<3�)�l�D>N`{�J@邟����f=����Sۂ��H"N<���'Ĵa�!��$�r(�[F΋�ڒǼ�>��_wq����šG��c[E.JR��W��׿q"��R�.��E([��$>�!&q��D`Y�|a|��~�'����+P��8�+GIEl?�s����U��l+;rSe{~�{�vI0X7�\i�vQ-�L������V��е��J\��Q�Iaw���	+��>t�&W�h��2�Y�R�^ e+x	�v��W��d�i�~����ܿ|Z��]��^iHܞ�!��O�馛��pH}���Pvk_p���%��#��`Q�Mo��zo
���O|�����%v�^N)ŝ�TS`sG���5X��p�#B�HvPp,J��'q��+K������]"q���>*�nr
g��:|���q���w�I
ք�>s�����^��������gW��r\�H�X�8D�렴v���y/�n��1m[�w(;�ت��Ӌ�.r�Ў���E����Қ`� M�-	3�J�1�pK.���y@q�ht�)�0�����;�7JBI2��XW׀��"7�f�a�<���y�u�}����r�A<�q������|����i��g-��/�)$q��;���S����$�-�rZ�@
�X@[g�O��x��{B�I�	\������V�Tѝ���Ѹ0��&&n�s������$e�z��b\r�{�w�����n}>�����un��%v�����n�짷c�;�\�$r�Ȕ�ɾҝ�����;���1�'�ΝJO���(�[����+^���2|7�jTA���%��3�E:�椞��<��I!�J\#\I���ϭ�C[>��F屢�k|t�_N$v�R�X�*a���m���P@H���WE�Pq�q�}���O��X�𠌄Cj$�b�K�P��.�8���ܧZn@g��Apȁ��9�q�9�H��4愡s�H�(�fC'����x�����ܖg�q�:t�7T���0E`�H��v�7u�A���?��^w����d.�-�~尌�|�̜1M��j��� ������bQ����Z�z��#q�_�ݩCM�|���йv_}-^�b5�(G�rFe�N$�Q7!u�*2ǧ�M2��G�V.Pg�����'�I��%Pus�eX?�&.6r�c�����9��<�:1=$��[��x��F��Ϭ�-�w(H\�8<���c��׹s�^c,q�t ��f�b�X;Ր�]s���ĉ;5+�ӏ�5�8�Sp���[�*���	3�:�*��ݿĺ�e�I�j��L�Ґ���9p�E`WHQ��@H���r!>��K����vղW��#�=�JT�{��N|泟�������n�_}X�c�$P���83!r��_&6d��P,q�_�Ć�%qz�I�@Ŷ6̿j.^�r5&w�`'��BّȨ�ʗ���b1�x��Ka%�zT�    IDAT�T��f�8��|w�� av1Q\��� 2�ĎX����c����Y'AwޅJR�n �2�H�*\�7�!s�ҽ�9V�؝[}궮�Y�f͚��+�������!<7I��7߼���� c����yG�IOb]
2x��k��.�M"'�~�hf˥	l�C���ذa�Te��4I"D�`L��}$���U�N�G�\w�!��$.�&�7��;��w�*Җ�?�W^y�,�\���-�я���|Aܯ���.��~����
]3�/���X�;�B��3���aD�츊�Mm���+q�kp��.X�ߵe����I��\L�g����S�F��9Bw��IQ#q6�����a(n�2W��Љx֏�jwj���`N�E�@�Ŗ�d��,m(�zk�t�1�\���}�Eo�k���x�K���Y�K��d�c ���Mzq�������������4�= � \b`$N��>��6��-JeYR��V�v�;�����zث�"�j�r��K�VQPF�Ll�1q�K������FBb��ާٿ/�#qLb�T.��/���"�#4��]�N֮��fM�Cn���1�T��$D��f|���睋@�"X��q|�曰��a1!)ႌc_,Vt���mP$p,�UG�.��Su�ҐH�p=�9.�R7�6o�����zS�+��C%1,2*�B���BF�Y1�9#�(���dA��$l~��I�X}CH\
�"��F�'����|�{6|֐�]T"[�oJ��.[����9iwn�ݵ�r�r���>��W\q�u������s3&��o��X,R�P��gw?�ۻ��e�x~��~\w�u=�A�$n(b�wO���@I\���!�tf����guJ%�^2�$	_����b'A�b�s�@%$.��jgM�N��MllQ���3$n`o�H:j{$��=q��+�]��!1�Eʬ�J]�6���.�8��e�<����Q�T��P@�ډ3�b����j\M�f�F�t��?~ �j�ˉV\Wk�8�3�H�$N�9����a�Usqꪗp��n�$��B�(�K�l�z@ţ ���˒��$�;�))!�l���T�8/�uL\���	-X�Z@�� �b����N�=&/���cO�?�I\6&͚5��W]uݩîP��N�oѢE��ַ�u�\���|>/A�{��֭l��=�쳥bCF<3���x� � �b`$N�Eֳ�}Үle���%�^u��/x2��ߴ%�$�.hk$���b�ɩ�v����!qd��P��%���=�J�4z߻����Dq9�1T6ڻ*p�@�c۳P���l%��UW�0q��n���/¦M]�-��� Y��d�m���S���j�����s�f�;��е�%��g?��ִ��@� e��X�5�"t:q��uv�#��3�^�]˪�e/�iӳE7O���������c�֌.�ܘGRM`�
�Q5�C�\#q����i۹3f�!��Ć���z�����#f�E�w�M7-)�˓�d0fV�-ӽ���.���3�p���j!�l;?��Ρ�$�8n���q���8]9XKL�8n�fj�L\�c٭�=$&�߽Eb䵈�!m;�t�{n��IB��+���N��˹����|�h�͜v��
�vE�B��jq^�����)��"�s,����>��|�6<�b5,�C5�Eέ�S�5���'q�]�^̘6�$N�%�X�}�KX�OWଗ��Ю2T�"�b$~ԇ���)��,0��+R�;U��N$dXʖ)K�!�-j�
xxL#�#���	�sY*���7�V��Jz*rl������/��ܩ��?���]w�uW���v���7��~���|��7��iI�
��E���y*C��T+�b駲���S����b[�e��{
�W	,�R��,+�R�eYT��K	���SN����|�@IgEB愸�b���d`$��j���z�B8h�I���z�6'*���Q�<��"���d}m��w�����9j_A`{$��TƧ����%�rY|����\��?.�?|i���Ȇ�l�<�^FKc��ɨl�mk߾������0J%.�bZ�ͳQ�QR<�-��\HC�"|a-�{mtԊ���N���]Ôa��Pn�����Ii�θQ�ݭ)=�Gȵ�H�<[�X�j
�b]��-��ƐTbx*��6��f��[9'{�w���#٩�����׿��/]1�KC��Wz�!o�ҥ'�J��(���� %���:M-�q,~ڶ��Y���m[�i*D�����g}k�g��S%=;�Rʱm���Y{iR�Ei��
��T�X�=����k��v:I�$I\}\� @�N1�$����Eҷ(='���cݻ#��:�cX�-{m��1Z�$���$qt�2��JR4i>�q�9��\-�~�<��|z�P')	���F�Q�M�u�L3c��^�?�߅���l���x��Ƭ&%aÙ�%�B>Q��^���^�����_��zee˂��M+M�ĥ���2DWJiQ��z�5��<P��{�S��x��
ZJY�J�4QpՖ hy�F�p���ׂ��nx����F�]d����ߎ��	܎�rֆO<�߾�կ~~G������f�[�l�����oy�{��6ZϗM�t	�����F���N�-J�M�+��zI�����$�NA��pa��qo���*��⃶5@ok���Ϫie���H��"��82V��8,�ƞ~ډ���BK��utu���u�����6�rrR�3�ܟ���;�/|>�O�d$�O>�߾�V<�̳"��Z+\�i���%qԷ�,��J�/����ז�7u���(o��e�^Xuc/M���\�I�I˶蒉-�"�ݡ��Z�Ҟ��N�-K)K%
*�-*�!�E,����%��I-U
�ᮢ����47���=ϱt�NX+IHxU�
�O6^�)w�]'3l�t�I_����%�]���~¢�K~|饗^�=�y����^ב��<�c٭l��Ic�C�4�c�h���\R*�#�2FN+���%8,�͠�����*:qR�1M0�Z�9������K�Y��$1w:G���j�ܨ2�5tfW&V,�}�������cT�I��%t�ή�:���������/eT;���-;'^޷Ԑ�XC[:H�]��}g���ZW����G��
�{�,���E[9	g�(�KU���-nڋ��KVO�f�����]�F��jI�Q��cu�d�����v���u��\���z�/��-�.��2-C}���������=#����v�l�+�dA�=8e8˳���m�sv$��]�6��R<�F�h}�L����_��� ����%�d�Į=��C��{��ʿ���!�m)p������� �bN8����\p@��و�7��]�{߯P�T`;t�값LBHǻ�}�1s�a�����/�B�ƫ7c��~�O~��ˆSU���~���W��;���8��U���C����o�ܜ�iK�����������S���|����p��۹�{��m,q{�a{�U�V��w�|��٧e/M��#.���N�58$�g>��p�T(�*�	_�M�,e[�̒iPH�&>V��/��T�hLY;���ׄ�)ƕI���,�a^����x�p��LM�x��0�	�v`Q���F�g�[n��Lpҷ��g�HY���D==Jb46�Q.w!JCQ�,��72��QY�$*0���W>,�EI1�������#%��h�5����I%�҉iG�{7t���hQ�:T~W2!�ٔ��]0l��+�RԲ.6]�i���2�Z�ײ��,3�0�	��R�,���$ ��B��۶Ei���}h�?�l��*��)��h��D��8�j�<H9��[�����!���_�UT�V;
�0F']u9.3��9��"�A��!)[�T��Q�,���x�ob`ZS�w����j-xSH��=��P���RM�R�~�lۜ�z9��Z�J˅�#Xv,�'�,��r��+Ea�����Jb�{��ތ́�$"\���gb�$��a{�V��+x��U*L=�0̛{��2+D��3,^r7J�**�B>� :q"i(���0~,���w���4��J�0n��-X�~l�E\[����u��V̜~.�䃘1�H�O��!�N嫢��6m؈�w�~��<���}�����477J)�8��ڥR�[�|������W���nݺ�*��$۶'�iڤI4�=]GU�+��\�?���y� �c�=��������n�r~C���^t�sϽp�=�.%�;y_#qY�z2�ַb��9�����}���T�.��ȹ�b�$?2)�AE�ԨH�:��]�O�'İ�K��,U�v*i�@T�b�eՌ
\�yN�	����)��y����~�5��-��/ -���2U#DW�$��y��H����bS�mn@cs����0�-쨢��)���V�*,���I�"�R!$/$Un��>��%.Q%8E/Gr�4`�����_0e�sj!7j� �0۱W+���KE��2r��$)Z�8�WkA�AZ#��_�v�RC$���Cz�nأ�E���R��Q$ЬC��T@��B�4�H�����ph_H8媐��0FT.�F(X� EZ."��Y*Y�2�k�d:��HR���&l)EpG�������&U��2��"�b'���FυU�$c�ﵻRE�QKe�J)��3�ϴm��`�$������Py>� (��S��~�ZVU�S^J��k]fZ��_��S��"���\(x2�Ϛ1��ehl�UlܰK���!���d֦���� �s�\F|g�~*���w���A���/�g?��Z�ZH �%54�Y�*�7�Z��ӏ��sfc��)p�9�$.����ڰ`���̛7�F��D��C=4aٲe���K$tǴ��^�V'�a8���Q�������������/�az����O�ǟ���wGl����۴|��������ϙ=��}���[�[��wEf��V�^�6I��x����Ľ1 �V�
�Hm�'�֜'�tX��|�,('El��r(8��D'P׹SŕWsˊU�.���*�I,*��B��nn���sZt3�"�C'������C��<�'��ۜ�E�)���n؊��_@��*]M�U�[&L��ԏM���:'g1�9E�V��oĩ�$T����&��OD��#?v<��Q�s�\ qP4������݉�R��5��]o�&�"9u,DaY��>�8�}��vh�J��h[J�-�\ "ZNm=Q�<��i׹�0q���St9�N���������o\#\Z�J1�ލ�k�нv-*�W�޲�INT�o[�I��nƠ:,ZB?�ǖ(Aw���#�Ǝ�7q
��aԘ���k��]]�\��ukQ^�����7�c�|
�_/f�3=Ӣn���$���:���YW)�Q�\�7�:e
��(�>�#Pf#��V���Ph�@�����u0u���"qYv*�ƴ:k����-8�(&'D�Xv����_x��v �o�	�t�<	�}X%1r�Z���#��3���,p�qtv�z��IZZh[$n��)Cn����ƍ�`��[�ͻ���#~�뮻
˖-kY�r��5k��y��� Z-���8vh����q����[K������Ňԅ:���B�6p��d?>�U�R۶�����̙3�p뭷n��7{e���?��_�����>ݐ���@&AЯ�.���}{H\�JL[�_��w��L2w�9�PO�G�SI��$��%�x),בt�Љ`��C�zp©���	G���н'R5���%��'tF)��[~�l����rF9G�q��CGj#�8	�|2F{0~0�	�96&���� /�A�c��߰�J!g��*v��+����R��y��W����!J��|K+�v8�L�{�$`�D��	�z�H�;(������m����>�MO>��}�8�KW��JKR��.�Z"��Q֜�li����,D��C�$����/U�?h2�9�=8b&�:AkX0�-����m$6�[=��?� *���+vaLc尌��R*�v�h��tD	*�F�e�4��9�YG�O���sG�}�ġ�(-k���E�m�����Q^#�j�ܛ~nE����Z�%��IH�T�bC6���/�=���$�������?��.(��MI��H�+c=
�2>3��$�ygV�X�X����R׸f��[MP�s�,����k����\��̞��@;��q$DN��5��3�,qC�N�g��y޼��ҝ:XSU���/XӧO��n�jO�4�������U.�� �j�*����J�R��}_ߦ(�T�PP������#��r�q㢳�>�o��`�� �ǐ�Ar��Fb�����sf��o�8������|e�@߀�Z�w6��!qzBeY�C��N�7~.�iK�h����� �F�X�P1F�uQ�t�UTƶb�;> ��s�$��?��	^JPП[�QO#H@�˱(�*�v36�b	6���hN��N�V�0y
Ɲy6�SOF���>?'O&R�S"�Y@6:����cX����^��@O��'�]�#1oĹ1q�D	�xH�yt�Bô#1���a4-+����SW��:)����cKݖ��# � �C�|[�y
[�-֬E>�`��1+J�D����(˦�H*���F:�o,r����D!�6���	8��1����&��dȳ���g��jU�퉇���������(��HH&m%J� ;��B#&�r28�t`�8���GwK��ă��}̴Dޏ�V>��'��7�CP�@3���.x5+(�*)��-#���Ȕ�5�-����1��K�b@L�����G��Ƿ�߰IZ�kA�p�1pK���
]�1qt�:ݣ,��.�E�&c�\���vm�CE�)��Y��]�}[J"�:����eK�J�H�2�z�\$خĜj��X'|8u$n��)�$�����;����Խ�7R�ӡh�!qC��0��ʕ+'�u��?�={�9��m�c����}=�zYL\?K�#��~�,JL\Ub�ΙЌ�$N�T^N!	LHp,U��6��q�8�]D�� ^`��ղ"eέ��q�!oG���Ƴ�ɿ��.Ʀ�݋QբL�nsڝ G���g��Py>"&2�z'~^m�d	؎#M^�у�K�܃Ⓩabރ])K�c�J�����I&(���2�N=α� �LE���6�ćOyC���>���������(:��� ��CX�翠s�ߡ*E4�@@�Z�	��Ӥ�Y�9�qO�h��t3R�>F�R���v���ޏƓ� Z'vq����G�T*Ǹ�+�t�1��>���橧0*N���HR��c�`��O�!o|p�!���x=���3л���kZU ��Vc�}�������^\�>��pZw��۸Ɓ-]x�u(��L�<�G��|����y����I�`�Zl�����#H�ݒd�0���P�7;u�$Ε�X5�6����Ť�,�=Jq���e1S$q�X���Ԋ�Ke�yL�4�=�z$�dKRP���|]�K.G��mD8jڑ����N$��ԅ�ؘ�a4%���7�lp�bŊ���;x�y�"�{��D���M�%��]'U�"�w�jI���)��Ter�.�.^j���F�c[q�����jEu�ZN��lt1X=��"D�݂$&�$C`K�.Y��_.��r	������u�`�;�L`��*kQZ�O�F����<Ua�܈.ؚ��}3��<����]�Q�8S0"Ij����=ޡ��i��w���c���b�䉎�R���O(�K,�b��P��Sv�F����$���z�Q���o.��.�i��X9�8U��d��Wњ��FMx�ܤt���b����Sq��/� i�鉕�f����cWb�O��P܂���/An�F40a�� �}l�T���#��.���IY����$S�G�%$Y�h�I6�b�M���W��ߟ���D+����B�Ԏ4�rp.rI������/�^��08�r��Y���OhjA� �ĥ�Qf�stu ����Y��c3�J!/���#qcB��d%S�C�>��A�&�#m�th1cf��K|g�3jIHE�ǾW�    IDAT�D�F,tQ,�Aޗ>"9�,��Y�U�P���p'q��-\�হs������l�C�{���=��K�{�?�=g�������7��O7�է�������(��@G�k����
ck#Yb	����Iu
[dAr��0IP,lni��s.è�N
'tʏ��'qS�1�I��6I,��&�tDb��mKc��Ũr�|3V��~�)�I�r�CrR,[��4�ѣ�|�޶Q�T�c|1c�zO�|Fw���.��ײ}(Ǒ��"�[��s�C�߬	\Y������D,"B��.��B�S�����Q:V�D2�$l#�iK�x5�ho^z	[�/B��*��l@���|�yfG[nХ!�@\uɑ"�$;:m��4�j`ʑH������qغ�MkP,u�i�h�&4��{g�cU�=�a���P}�)4��E	��BwK+��ۑ?�|`�xĎ�jZE��$Λ���v�E4�Z�L: د��!���tkT�����_�C��$TUH%S��?ݞBB�BZd�f|X��Ǿ�}��$n �P�b!>��Eщ��������x�(01c7�8Z�H�(1"^t��,�I�$c3{&�H��]�L&�	�?�����l�A��@jrXӐ|wٜ٘1m�ݩ�1q�-�᪫���n�2��������Y������gϞ-b���+��]'N,&\e����ț��*����"6"�!.R����>^�J ��8:~-��Q�+�-K\;ΙЂ��N\&�P�q0-x0[6�6P�o"~�l4�q&�Gi�݊�.t>����c\���Z�Z��B�"��B�ME@��M�-ÖgA3e$*.:[[1��I6ݴ�&S7�r�o���ǰ��5���g���I�#݄T9p��j5V�໰_Z�ִ�JgT�A�B�����`c�ื���g�ր�b����d
a\��{ /?�����J�O�ЈIS�c�ѳ�C� �9$��(G�^T��vo�,���#:�^F��82���j@�Z��#�Օ��j���F�r�ѳp��?4�P�-��'�����oX��_�v�X�D�=e*&����aG"�|�v�"������Xv��[�h�(V4L?
>�`�LT�&PD�N�ha,�O�_܃d��b�S@��1�ܓ�s�Qe�������6�������C�7��P�{�Cɷ$��KC�f�Y���X�2g}�����$�8&1,q�R��NC�ԍu?�)�<�'�[���֫�vr���wgG�Z_Y�!���L��o�`�f�vt���LF%+��+L���5��:!k�����a&]?�Z�P�N�es.v$n���ϛwհ����ھt=C�����ƽ������.�=����Z�2_~C	Y�{:�3�umY�ә����dc�9#g��aPT��_�NUi�ƴ���^GK���B&��@~�d���i'�0��_��O�A�qk9!�dU�V��;�b�O�I�H�%�u�RJ�#���c#�CIr�J�(8�����O��	��(�ĉ�;J�R���+��7n��~=���l�(�.>�4L|�y���<������|�v��m��(�!��C1�0s&�������	aj��V�y׮Ú��ol|�ɂ��T\�l�GD�\Zc���fD��1���O��� "_^��������h�J��yZ\��n�(8MB�c�*%�h��j5�9'���!j��O=�[�
�4�X��
����g���?�ڴK?Y
���0
�\����N�e1�ڴR����x��o�Pڊ�려<p��h|�;���%�e������7����C����F�����0���IG!�D>�����w/��E�0:,��sl�R��EٷD��M4�c����<�\�&�������VJ�ɋŒ�d�$��Ò��>���w�J7u���k;#��$N��$��F�OV9c��8��0�IܿΛw��}|J��nߐ�}���ް!q۶�enU)Ek]7q� ��sltvR薖8)e5�X��j*��F#�#az5wք\��NՖ��c,NU�T�
�-$�%��dP7��g6���a�wM�$���?�)��?�f�MbP`���	�F�`{�|G,t��T�5�0��>���IH�܏Kw���[nE��M��N���Q��3���M@sV�y?ʛ6��%��N��-[�p�<*��x�~���7�9��0q�R,�&)
�PO?���X���g1�I��cyaR��V��!2� B����5�	�.�]p!�l){O��N$[^B�v#P."E\U�� �R@"�r."�Z+�EG+Z�
p����9�.��q�E���?��Uk�%!��?�$.60���0�ҏ-�R'e��}��kK�t��܊��ȶ�P�'Y��:�i�|���vLb��8�BTb��Zr�������$��h�M�F��ߟ���e��o��&��/"�!��D�,"Ȗ'���W��<tWc4��,q�\��٫�3Z��X�/��{q5�JQ�CtV�~�2U�7�'�*����N�o��Y��s}-k���-��#��S�Ag���4Z���,q�s��Ծ#�0o�U���S�>w����s]nH���K�yk�@wj}}H�b�v�ihjl��?�M��R����e�S�rH� �r��RD!�o�č	i�k�$���Sl�$��u����BGw(�q�q������>��Q&�sE`��x�{?@�'�����z�l��B\��,�F5*���|�%�\lln��_�6�!*�B�RA�x�7��_�D+���$ᢛ�R�B9BC����&$v�F�F�*8�4P�
h}�	}�ہ&�{
Tq:6k��w7|���0�3m���P�V�z�RH�p&>0�U*��dWPl�c}�ǡ'��N?�3����_!�n���s��Yu<�B�W=X�-.Z�K���"���)�����v�G)��T9�-[ќ(xJ(I�+�][�N:G|�����lf�?��v��*�$��t&L��7��i۴��F뺗Q`�$����6[6�n
��8�O�
9WN�Nx�����и~
v(�!�>�b���᧑����͘�I��Y�e���KU4(mhG���q��j�H�����N<�d>���(Ԉ/I[�^�S'��6�?�����-q�r^_A�ם�큽O�າy}����Yk�5� ZZy�,�5gN-;u����Λ;�ʯ��S�>w����s]nH܎�����D��x?.z�;���?���^|�%T���~a�J)��t�@,^����O��H�N�C���f*��SG��-0;E�&�&1��P?�\4.u���NnE`�KX������Sh�	ʊe�<��W{)���$�d�#k��mt67��O\
�r:Isc`!B#'�?']O<�_�V��Y��#b��������tu#O�\lɹ�G�`ڻ���o@� `�t��E���-����[1*g�T���>|8���ƼN��Sԕںb�A��r�ȏ��$�Q^׆ f�E;�B�e��K_t���-d�%�d�"�
%NH�r�X�� ���s5��HUEȘ�A%�~�z��jA�C�Ao�?�O9MRXKqU��Ng;*�~����n$A�c�ńw��|J�F8�u��sO�/_�DEإ8� U��*�
M����u�X��]�����Xy�7�V.�wKf���������J����(��º������0�*lx�	�}a�=�L���eU��/��G��5�׮�h����r�3FŢli���lw��eqmٹ_���7>.�����ڨ�$N�=#�/	r�g���Mg�Z熏%����]�o�����ݾ!q�\���a�N����Lbö'�\ࡽ}+�?�l���o�a�OƸ1X��>� ���xy��]R����D��G��[K��v*q�h�N\؎s�kƅ9��J�XH�$a�6%�i(����,������A�����ݯ/?���駑��/���z<��P�]�L+%�4�Z��(S�t�t|�%�A�4�T�(R�u�:l��n�}�A�:;�v�O
��b�)TOHm��S��l<��L��p���X><ۇS�{n+���ۨ��Q�o)���`�	<f��PB�!�*q#3��Y�l3���	6��Kp��Ȥ�(��p��H7��Ģʯ��"f�bj#����O�S�z�l��2~Q�=kA��h(�C�>z�T�Sn�j҉� vs���?�x��;hlD�:V7@x�	���;>��j��	ͧ����z����5��J�T��g<����2y�%<<t�pstsF��][.����	x���k�վ?�1��$�Vx*A.	$6��U��3(�}�A8�sW E9�$B�ֺ����=�b�����s�C��St)5�@V˨���G?@�~��jf��Ɉ��b�L�R���%\�����y��+D�px������%�(Il�)�5�H����?{��s�}�����7$n���7,:q����ٳ�o^9	�t��{�onl�I�?�}��]lnnF{w����?�	_��P�+4��Wӳ�P#q��o�K�Z�X%���'�M}a)�^*%�$�vP�R�N%�k:�|��fiBiG�{��uR�A�O�@�C7��;(%e�q���
:�]�����,��J�B�
p�������?{�fUyn�v��ieh�-�b�5��ƨ1�^���n�MSј���o�1�FM��5�h쨀� m�L?e��Y���`,�`8��30�s���.��ֻ޵r5C9Jш���zV��,V>�O��I�V�}���t	�?�W�Űi�h��#оr��@�!�*)=�eX:/��jT�lF�N�Z��3	�	�#���"�l�=x���/#VA��Ѓ@t	��v�f�#N#�8�)CDC^#bJC�!Lڋ�pX�W�9��m  ��-)i����A��P��8vC_��o 0p�T���%[�k} M�<��R?@)_@�A���3�m@��I����s���7A��c��ǭ�T*X[�1���PԱJ��!]�"0�N�{�>xZ;,��-8�J� #���Pw��0ⴳ��$��6��23���2F�w ��rP]�F�1�#@��t̽��mo����2�&r��1�d'M@=�����o°�7��*݁z�3q�A��c��Ira�&M��'^���)���𷁸�S��/\�p��S���{�z ���t����DL�K4"������ڟluNХ �r]'�i&�;��*�َ��\��A6���;���p�i�b�FJ<OK{Ӧ��g�|s澅��x�ZU	� Nldٝ�2q�7���^LK�Fd��^���$��޽��mw�y���@�w��}�O���cɔ&^�H%E&�}�"`�*t<�V��	T�E�ˈ"N��ǈ/	�3`��R����u(?��?�O��5�V\-`׍lx� ��:tva�l4[:�{4�r:� %F4'Q��Ϙ{��h�b8]]0#������C�'0K:h���Y!@�Z���>u�b�z� 9S����2l��E��<4i�N�`Y��6��&�8K%4���@��Q6��3iC�!��+��0۝u6���@T��3���Q�Qe��[m�t<�=��V��Ӭ��������Q�H
�(��8�]� ��v,~�Xv	z�nXUN�b�;�"q5��!�=	�cƪ��$Sv���{�$Z���B��-;]���4�*Tc��^�8V��r\�2����G�ڤ;%�l�^����S��;0�JE�q�|s.�j�W *e! f�Q,~n�4�������^���_c�ީ��_5q��p��8If��^[o���Aʩ�ĩ�&DqZL����w��!+�n�L�]_�8��>��ﶍ~l#��}lC�elxNc�G��w��ם�ʵ-�1i�I��Z�mW�������'�Ho���10���5���J��cĈ��m�.���q�~{>jk��Pp��R��3p߃b���%���?.�T'�ʩ ����R��@���s�˯��IO"���z�9(������^��_b�8/��=�s����~0A�2*::�z�d�{�	���%�V�%I��ƍ�Nǝs�@���J�_W��֮v`�L,��*K�ֻ��]��:B� ��/ԠR�P���v'������|_p��J�Y�:�p�U�f���T�KdW�je�\s,S�_�0'
��R�2��d2Cb��i��QB&�qr�����C��Cb��N�J�H�Y	Qg���2
�����TI]��8��Ul��H�.��G@紗PSlCވ�z�sX��q֙�{<`�k��P�*����C�O�6a�g eq�k�)�IhDh.�(zFw0h{��A��<�f�q+
I'b�f�
^��>��JŇo����|�[H���+z���v�b����(͚W��R�a�/^ �%U�J�96��Yyx
f����V��2�i:m�@-a���V���43\i�,�yV�̺S�^٩:JdS���@��/��^=�nfX�=ʒd�gSo�ÑӒl���3�6C�߳~v*�8�B�L\vt���ɤɓ�|�e�ݼ%<����G7�@�G7�[�,X0f��~���H?m�	�e�R� .=y�nG�1 N]���~�Zuu\���1����{b�]�a�N;��7�����3gV4�D����Ԟ�c��a�n��2�G���J&.q�2;��0������w2�AV�)�`z ;��0�s�#��S'�D���oE��&P�ݐ:�z��X}�}X��aL}TAL�CG{��\Us��=�T`�]�B5��� L�e��o��ڧ�Yϡ�lTW
��ʡ����Lh8�󰏜 �J�>����W|�⅒"a�	
����`h�0���EB�F
�	���U�����+�5n����	����6�q4sa�����vFr	Hd˂���-j	�Ǖ qtDCFc����g?��a�R���8�ǧi��|3_�꙯�K����䡣���<���	�����E4���_}}�.Xq��S�D���B4��:�>s20xL���A+������*�[P&�s_)K�H�S��N8�q'"��AD��~�Z���1��?�Y�
�����Ps��v܉���rJ�r1^�ߟ�X���@���g�q-�IE�a	�x��8���Tى�H�L���]@\������r�f�,�N]YU=����V .�"�F�=�]�\.c�g��������onn�Rw��8޶�lq�Po��7o�ةO���矻˅�K�fJ'�D��z(*���}�@���h��,�ħ���{6ƍ���"-�K/MC�F̝���"�|;��q��������Ɔ�� �<���#��A���%�B�p�e�P*�qRZ%�[�
���'GxI ��t݆ϮR�A��c��{�jk��:|�-�Tz3~盯c�S�b��W�3�b,�8.�ȡ�o=�~
j�8�s�F��҅7/�&�V4���9��Bj�T�{�P>n�}! %��K,,���l1�/�N�
��RK��e�+�*Y�����m�������e��*�Φۖĉ᧜�3�Ӂ%�Ey�tx�׀b+¥����>f�jA��:8�l4�!ش���$���"�5���ʱ#�a��1��ߵ��>�!ǟ
��i`2��ix��ѿ���@�rP���������D80���o�������38c��r���:G�]c;�D�`�q��tۍhz��	J�L���%��bO�k\5��N�֦�88A��k�ޞذ�D�]EH����V�I�'}��.��̩v���6�نv����󗌛����/<�ܽߩ�!!��iͺ'�w����c���'n=&�7���JC������p�Ab�x��٘;g6�-[�r���V�ឆ�:j����(ӥ����ĩr����Ā��Ȇ0qG &}�M0QJt=^���Xs\J�|��p�    IDAT%j$�F�N��W�{�q,�A�+%I���i(��;�����(A��qp�������Ps��	�~cE��W?4M�^E����h#���}O9	GD.`ے�u�b�.��d)b[Gxp	֘�9٤P1r�N�KR$��1+��B�)`G�pnO/]��̽AK�R�����ℽS̎����2��D2:!�_Mq]=F|0��N@��@�>�����@�j�yI1vY#�Ly ˞~
����������q�9c	Y��E,��/��yV�KʲFL���$��Z\u���;<���e��r/Oô���J	&u�9?�m�f٨?�04�t��U�&��N`�b,��-�Z5fL�b������Ϝ㘣���il8���6`�tL��w�-�A�Jpi	C��������N�A{����cu�36.{�o%�N]V.��0qޤɓ�����Q�;�������|�{0wѢ�L}���?o� ��>���S��75��X� ��&��w�N�f��y8����6���֭mFWW��*�}�a|?
($�=��&�wqm`b-F6�BM�%�{�7�Z��O>o�8~GlK4����켌����;��Q��9�*�`c}�L]��p� l��Q��ӆ�����w�e8�4�.`q#����-B] �T�86Zj��p���=�XJ{�b�~q-�����0�4fsA"�?�&�ءLϲ��t�Y���Z1��R%W�YKE�)�#�r)@#���;�����9�C�Z �@Dgt��f��!}�%ǀӧ� i��1;b�����#�B�j0<��
�W_��)�Bo���8�г/Bñ'�X+A�y����/�>nP��Nۈ��"���ֹ9���|�La=�ٲ!�Ax����bpكY.����#hV:��Ŏ_<��.1lh<��2J��Ǣ<��kA�N����@��]1��S�����80}fԶb��A�7P{�+%��%KVU��Y�R��9R����$'g+q=��k�z����"
aB@\e����y�e?���8޶�lq�Po���ظ��)�q�y�W�Oq�H���Ygf��F������07������т����8����[~�����X�e9��|�a�:_��RE�g�d�2��6M\o��nl�(&� �.�d!X�\����ߜ��#G(a�-Bl)�؁��	��\%B�P8RqRJ���^���\�0Alh��C��{c�A�;��B6~І��#%���x�1�+���(�!:���p�It��E�q��^:��#���1�<���H��#)�	;�+�"l�4-PQES�H�3A��QJ(���ɽ�����	Ӗ�tJ*b{�eN�t���P���J>�CL���텍?�?ӂ�%�<:��C0l���p��@�~�3T��h[�����A�[q�������FZ�x�+X�������/ Nű�&�H��Q��AG~>{2пe��Z7,�MŌ?ގ~]
Q����6�c5{_<28�)�\�K�}-����%��>\k���uv���u�D��xq�@�G��n� v���/(�6-�ĮХ����+ҝ-K��j��i�ֳY1�~�VOÃz�r�ذ�O�V]N-O�k�W\�������6����6���������1塩8��/��SN%����-�z����r�V⤃��ӽ����vL88v�18��3в���z3fNMLeuÖ�)Ӷ��꘮�:2q�� ��D��8�a��b䰁�
�XN�!���P�u��p����-�a�p�@��jf,������"�$@��5)+��"��E�cb�B�b��r`�U(i�
u|���������]h$0����Ͽ�:�Ͽ��I�r� �p��u�@�`����M����+�݆�5-�C8���J���#�=6`�F��d�'��jN �!�S`N�e�C ��S8%���Y4r�ȝ�ta�Z�T�.->Z�T��PKg9�+h"��q���B-�P�Z? ���C݄���Z�K%@��930�����;�x4{"PW��d�i�؎�'a�Ï�&*ID�,:Ҳa�rjA��j����/*���`����+��� E�E�[��?w
l�Ek9���`�T�^�J�`�.�$�5��"i��1�::�qZ�,�������%hț��K2>v�=20$-z����BtA�x�	�������^.t��z��n� �ɓ��x�eWo9�˶=�(F`��(Fy����������:���v��La���e�Fp"�OO�����~[D{��1q���5i�:�:�H�y֩>x�(D�Qݑ��z}⊸�?����ʹ�COH��
��*�@5	�/����G4�M���2m%�t�Y�ch��b�4򑳔n��|'l�b�t�$�%Ǩ�^��Dw��UhqL>p?=�$��@ ����@+w��`��:��,,�}${O=1Vt|�.	�J͘v����`	�{Lh�Ć��|��ȁ�)��X��u������̞�%�K�p�y���qc7d7��)�:�)���bP�����,T#"i��X>1�2��Z�[�8�RE��ˆ��hA�p�(�~��@�� 
�§,����͍�0��c0䳟��A`��F���(��;�b����Ӱ�;E��m5����K_��ߧW�
Г���f���&���S�5D�
�\�ul41��y>0n7D9. �)sD�C ��d��")
�H*4�B��ɢ�P$��S���ehh
V>�0�eT���	[b�Bo9��DG�8r���)L\O�JƤ���w����瑬���#ik��-�;uMssi���?�x�~�O7�vm3��6�uk��Eo�������E}u\L[Pv(:&���Y"��DGՒz��K�D�>|"@��]�YY��q������g���5U��g��8v�D�m-���߁G�>� K�d�XDڌL\b�%S�eW�%Xp�u���E�h)�{�6<�a�!\T�f�qP�e��<�D/�����	|#�AF��ySC��g���C[���1��#Pw��@}�t�
w�W�w���K.����H�.�\��;�|�E���Z6ִZ�|�^s����.hq���@+0a'��I�k	�7˷�)�KVm;MnN�Jb��PES�d����F5�IJk'@�,��Ĝ��L��5��U��G�h�`�U|_����%/<�>��2SKE�9X��.a�thv����Ջ��b0��jEhM˱�/ż�_ň����c�F�X�$��͹x��]��A'
V����k��D^��+�v��%�?�/|�����/Í�h��OPzu��!�z���:T���t��0��ây�G�G���E�����K=K���6d����UOJ�A#,�_��_^+	$��!�|��������O�4Wi�-��z��]]����u�89x��1�1�E	_���K�C��~�ܼ�xפ;�w���~�5�?��u�G`���1ܪ�a���v�w�C:����A�9s?�:'��r�O�
A��FѰ���85�*F��~m*�� ��MQ�cP�@��[C�uc�a �$3��(M�h��[dhЙ"0"js�Sl�)LNf˗`�7"|k
V�dSCY%��ѪŪ"��0�D&Qj��8?2Qa�Md��Ð]Fc��O�_��C:5�(�������>u���_���^@䈗0����uX{�������>Zj�`�Q0��NC��v�Y�܎��-/��y%����I1��P�T��ބ �lJZ��5�m�EK�ݸ�����4��[/OC���:˼>L#�<�1h�&3k�t,�jp�����ٍL?5�E��
#�}	0p��q����`�nCشF�Wl5�h,{���4����ޗ�u7�.P$��h��+f͆3zƜp��nH�����ʞX�������敨3}T�2��G9 49�Gb�/~	5�U)��v�����a/X����@��<d�p�:��+�j�ݗނ�1gS�!�qdU�[�ISƨ�T�:�t15�ln�G��%h��vt��*�V �>�K�x��8��!��8�g�g>��r���T6��ݤu�O�&�2м�?) n�]�����K'~�O�m��hG`��h�{��ڲ��y��n8�ܯ��y��.�'Q�1��A/��V'b�J��QD[3�S�oeL���xd%u�R������Ga��X��	o�zK�A%j�l�^�C)�Qg[��L�4�5��_���4b������W|�q,�?�GE�����50+f�C���ƺ�"ꝁ�Z��`���v�x�
��;����ѧ�}����Bʺ�U�����_G�� ���@�|�*���:t��j:��"S�Ît�����TI)�Z�<� �W������nkF!�Qc�<� &�j�ݍ07>Oi]���S{���1��G �b�c�ĺ�3Q�щ�^��3�a��0	��L���M)3Z�z��U[�q��*�� ��aZ ��Ɗ{�Ĳ�������$��_�B5*���PCy�p�qե�9���|d������|��к���}0��S�}�E̼U�0R.b����5 }�N�tx�LƚlW�`�1�A�〾��u�^@�\L��0��9OGb�hqt�����s�Fm/�R�c8�eJ�4��FΎ+̰8���*$��4� V�.q���l�;^�������i�(�g�!�ä��Jod�#H	{#�~��b,Z"&�qy7'��l�F����33�5�O�T��64�6걡ٺʩ)�'^v�7�lۡ�:	�K�=�C�˶:Ux3�t[��ճ�D���+�Jۇ��e��� ���M��_f��w��d��ｷ�!��Ͻ�3��g�?{���x�g�}�~�1�Y�X������{�"I$W���������QNי ��(N��4�v�+m�{��Ͻ�['Dz5�H������6�.4C��j�I���J+��6��{o�r����[F���9�r������oş�r�>f.Y�ٳ�H��f٢���w���,F$vKЌ����;��hs6r^$��FJ1� a'i�ÌuTi1B������^��;	' ÆR�T�ȿ�����s(�QcP�Ct�r�����΂1|$��Z:qE<־�'^���+a�:�s\�����s��x��@�vbRLʁY�֠���u�T�6�ܴ5n�O��n
KV�c����<���������UrBo.ĊG��ʬ7a�� ��χf�F��E��"f�zl�P��eMOװ�������!�#v�Q"��ȳQ��i�y�$hs�B_j�h�Ak�D{�4C;5'��i"���
�]���X���"X��{�v
p������u�f����[nD�89��<#q�Ib�0�|�i���@./��Z[Q|�I̹��ȅ&J����=�H�|�Di��<M#���t!�ukaq�⊊g˱<��x�ׄ��{�����n ��TQ����1�o@�l�vP�-��8����m7��IT�=Qے�i���,�N��
G�F ?��Q�q�?�T��M���/���oۃ�r6;�[7�w*m�cG�m�q�錚7N|�ub�Dj���Pm$����7�����@�[�t�wr�=���]�����5kRz��]�����;|b=J'۷��^��c�З�A�ʎ74M�>Ո�H��ӟT|655���1���8�h��������k.���'��h6	��}��sR]�� � O�߆�f|�ƃ86kd��H2&�e2�/a��a���ᘣĒ%�1rx�㯘���q�M7��9o��_��ͭp���e�	]rL�+vk|�:08ٲ�`�
4N{M�aT82�^o���*�+_*�}��M��P���pڹ�0�7��mŠ}�/��k�zk�ςS
��&�aC0�}��Ч?��Gƀ��K��e1�̑h��]:l��1򨣡�i�����w��}䤺|)�f�B�����mE�Uʾ %ݱ�T���Q�#v��ΌsP�=�Gq9�����X1�n�K� ��PE��F]3Y��-�BX�,�j�X�����C1�s��F����r�N�*tN�_|��Z;�2��a��=����@Gࣆ�0&"�5����Xt��ȗ*�D�!��S?l7�]����q�]�/��Ƨ���s�>r�T�~{�� jjC��v��mx��k`Ν��b9�Ekl 9cO?�{<"�E��TDV{޼�ft�9n�/���c�y5u���ã��u��.vs(Vp�׾-��48�i�-��G������63��uۧ Nil�8��c��B�$�Wo>ܨݣ�_�'z8&|H�����*K��{eI�q�e��wM�|�ĉ?��f|�~�_����]�|��e˖/����iq�A�q��t8E%�Ɨ�~i{r��%t��;C�Y]׍$'Ɏ�0�v�4W>�^x᪏| 6`��ĵθ�?�kf^nW��]�c��X�K08�7�nl�P|2��N�B>� ����u��V���4)~��W��(3��i�G�E3Bۆ� �%��(K��+�Տ���A�K���ą,���q�	��Yg���U��������ǔ)Sp����\˱p�o��?�$C��q|d�+;� �Z1j�T,�)�������"��	�N��&O>�%ݍ*��`�I�@�ԧ���-W� �d ��[�E�Q^�L�=r#����#�<eAAV����?�y�V*p�d�i�)�|Á;f�`p��2T�<����������Ytv!���Sǅַ�  	f^�ig�te��@[+��	M�����48�.�>�z8Z��~H����p"�� m��� �u���q{�bWHa>˖~	X�����	q������@1�?HB�e��F!"�9�c��w#�=�A?�Q��;�s���H�+/&'.�U��ޘ�u��	H6�<�G����� 3O�����B˖
0�<���ѯԅ�XG�]@n�0�Ӏ�z�&���8��1��k�EQ��x�s.P�݌jfb����ˑhW�:����Î��?�`��ѱ]/?���#����e(�X����Y̙<3�]�ƚ�Jc��G��N�~��R�_��W*tt�r�j4�Z��>��|���O��&�5��/����x��`ٲe�U�Vjll�`���K�.�w�ҥ;���&��u��4UM_�u˶m��}��!u6n���� J�m��k��~}�u��������6;z*θjb����ye8���]��Zߗ��9��oy?�� E�Uf���5wE����^ud`ԡ��}"ۖT�I`��8Y�j��8Y��	q)����c���r�����q�Y��_�t7^x៸��S�N���W|�ۗ`���=����Y�s]xq�%��q4��s`��$Hq�M���Dm��ER� 'Y����lB�}�<�,������ag�4B{����~��Q8�{y�J��Y��9W�cX�o�x=�7�@� �C4K-[΂O_?@`�Q7vw>�(`��
0	�����"[�Y拕��j|����.=��\B�R�4X�klD��Ϡm�4$���U:�j�Fu�:�pB��F�2˂N,�ęeTL�]�?摟���S��Kl�U�˱�O��/I\�U��f U��s�2}�{V{�(�i8h�,��#�:
���t~/[�= ��T%ȱ��Jy�G�a�@�*���X��+E�8D԰~�s�9�a,�C���Y�����`��!׶UZ�0�E��xl3���p9��4��Xu���r�0�{���$���!*�s����y�@���ۙ6/�nQ	%��}�) .|IR����?/�XZ�8t��ACG{��X�����s/��7羅J9�[�����D0q�]w�u���/���4�͟?�fɒ%#�.]:���q�~jݺu���rmE}�a��X�.D���6f.���j��s���w�m�_�򗿼�d߇��M�`�Jj    IDAT���^���U�����<d�@��iv��?f8�~f#��?�bW�����JZ�n����Ҩt�W��36��C!}�L�m
�W�Ì���%���A���]����جIC�d7��|�����;����hl��^u��>���;p��+pС����7��6�Z���
;���hL< �������8��G�4vK�G����1,���LP]l1J0�3�r"���NU�'.���`U�Y�x��݅�C��a������Tԅ�nV�q�;��P� �f����"�N�T����Y
��Z�����S�EMg���H,�ʡ��\�0Dk%��}�G���P��^��W�-n���N߃�NCi���ɕ�6�u8z��0j��h'A�Z��1˟ym�/w�	K0�@�Q�����#�& �5TLf3h�e�$�   H�h��w�ٰ;F�.m��j��Ɣ�h޳����1r;I	>K�օO��<���5�=f`0��D�u���b��0`�g�wO�6Oo9�kʪ&�� ;d5e��k*����J��G��%������T�eǅ���}���;
�J�	��������a-���6�9�>�����k���N�q�4��VW�Ѵ��ī����x�݉au���wb�cO��\�(5Ϥ1���U��|n(�D�f�41'41����P"�6�AT^���9�B�^y�4)��q�/�/:]�4gY!�S}��px� ^�>wM�Ͻ�*:�J��u�8�f�mn
'O�Ӕ�.��ɛ

>��/\�J���SN����Bi&��J�angg�H�J����q<��my^R�ɲxu�$�#�c���a3QV��}~'���wq������{�5�|SS�-��A\y���z�^�)�<����i�(<�ax�p����n���������z=f����F��?�����V��$J��
'f�F%:z��pB9�+=˖�����T�O�+�]�e��ꎹ���c��ej8��'��������b��������w
{�	\�����A��7a�=��
��
a�2PfÃFۃP�%�z]��k�WnW�\�����5-6b���ď�׫�q�U���8�0qy��&�Ry�Lz,���Ig�:)��v,��.��<��r	~��CC��/Fr0�zЯ?`�+FF�ݭi݂��&�atΨ�k��O`�3��hjBm�� ��k��F�N`��e5t�8r���>�'�� ����A�`vSI��p�4+#�N�!��OA�,_��W_��צ#\��Jr�3�󆌏�en�}f���_��Dp�B1�	ǭƪ��p��x���W#1�3vŮ���$~�j;�g&�2������,�z�	�����(pr�l�-y��p �xЯA�-�˞fe?h����A�ٺ5�|�%,z�	8����}O��&��~q���w�	@]�؄x�"�|�/>��oĀ�V~�D ���3�`��#Qr����q�[��O��_�&<�d�&�,�>s��78+V���)*a���:lɂB#R�e	�x)�Z�/\p���3�1t+}�93Q��-�B��g��^w/_A���y�GȜu���.� 4®cw�E^�]v�^̤y�di76S��gzf��0��͋����������W�V�Y<q��bzޤfx�T�X�(�-�n����=|P�N(�~���oy��N��{���S���l�TM��jl��>�y����tt��-�j@k9@�Mݲ�(��m��l��C"�(�c��>7��'?���%��x�'�UY=�$�@�Tt��2C�P6/�4!z�z�[>��~����E�f��ፕ1�pɏ�Ey����[��JPf\���
ĩ"��	S.�4��Kio�1o�#���Ndv^8&t�vW$������{��_�������a�.;`�ko����x�噸���b�[KD|��]����Q��I��xh(w�Ё58����V�&O:г씁8���#��g�3��ׯ/Ɯ�`�� � �{�gl�f۴����&-K�"Zۊ��C�c��ԅ�6)���(Bԧ#������~�8���p�s�w
��,Q�.º�_�ʗ_ �'P ��X%��F������b�ڪ����Q#0x���v�I�y�Tɔ���!P�t�rn!H
�K�5g>ֽ�ʍ��׬F��
ҭ饙��΂�.�b\�	���JtHSH��c��T�a�գl�P�ʣ~�]1�� cFn�����t��3�r	�3M3g����D�Gߺ=��4Qp�:���z��C1x�=Ѱ��b ,��v<��$�<*%ifi�E4>�,��GpİXG�v����8H�IJ-�X|�dT�|��bw�J��Kr�bD���~�i���_�0��-�!�6�����<���?�BHG��w�i�	�y]$�xn<��e�u��g��P�;��`^~�e1�>��1n���b�G)�q۟&�w�-�*��m� N�bD�v�\L��㗾���s���Fc$K��W≧��F&S�e9' NCl�����S#Әe?����/#c�e/��x�{�Ĉ(+�5AR_;{v�����o��g�v�-xͳd������{�o�w)�e�������?��v�j�ނ^���[���kߺ�B��@Vѩ�hA� ��x���+��4q=�m����ת�����%�8�[W"���&"v��W��gS��6��S8��?���,���n���B�`a� ȹ�[�1n���/�N;� �Q�A���sq������G����J%��⨲ �La�.�f�a�E �4,�[(Z6�}ǍE��!�#2L��~>뮕�� �Sm:u:�2�^����#hZ�*���bua���#TU�����Ѩ5
=��W�8��c�A3Z_���eKо|1�6TӮ��D
��&�'�n�s�'�k��tz�,ru}�� w@�G��6|8з KUH-/hcѲX�h�@��Ft�Y���&$p}n��ioK���p���\�,/ҌU��R���Z�A,PlpV*Fdm��5��7�Ϩ�1�q ���?)�� ^��+V�e�Bxk�@��K�@'��4��1ĚC'#�Y����A��E���(����8����`�);oW4+Wc��׬BԹn��
�H"v�k,IM_��#����0�!��bb��iȵ5˘e�타8>��������G��?V�c�]%�͝���S&��K6��oF�	��?G-�p�·�*�ԃ7�z���U�~|Օ3F9:��3�)�������ĥ�#�Q�eժgߖ���6�
֮��Iw^���_��n,�N�ī]4��D���V�^0ac��8��#Z-�(J�J�����6~���&#��|E(�K�n���`��$��o�������9���[��d�#��y�OQ����iJ�W�嗯�e��aSN��~��(l=�U������1�ܯ�b�sꄙ�Ê 	��x㫲��3&n�q��LC2%>R���O)� �Z��hGΦI����c�]�a�w@UU���ޜ7K�4��u!M]�#�t!"��}A˩�g)�cM��c/��Ȍ�+�t�:�P��V7TF(�ϔ��,a���ż9�$�^c<�9�W��J�UyF91�=FU�FJ4�J�Jy�����Pa(Y�T������T�z�Y1,�a�wF�5�E ��qj�z��*[���KPeHs�����6��+�����A��(?��3�+���)�TX2\�٢�|g&l�f�*�dw�	#F��Ϧ�%}�$N���S =c��d݂�����ƶa�ס�:i��9d�Ȟ�������E,z`2�aXaO�p�貙Ok�8�K�DM�s�Zm5P�!�T�1���qŇ�U���áE��I�GBG�t�օ��n� �L�n��o*r6�W�0d���{{�� ��݆G�]�9WE�>
�f�u|I'l(��(@��<�S��/�B|ἳ徣�r�C���nº浨���o|'��Yw�@>�,~�ӫ���]��2q��,��uͳ0i�wڿ����1���(`T��<K*�,,��ݤ�4��!���*:S����a�9�n�y:�xG�I?���kR�&�c�ɦ�6Ľ���d��c����^�oYN����\���g�R�&�+�����Z*�5���0�	W��1q�v��"�L,��3l���_����-eR��D�B�K2D���v(5�ܪ�8C��ӔH���)抍7a��� ��p;ﰽ��[׵��W_��QD�vXӲ��0�UN������� G�@nB#�!����2f����-ѦU"	�E��L*⋕�m��,b��)����4
���Ŏ�X@�I�* ��`�pT$����
��(8�uXa�ZZ��!¸�$
I��"Jc��$�]"�R�-C�E�N �'H��Άa��t%��[>��b�G���Yk��`��d�t�eK"ɹ�H���/c�2��2�L�K1td��$la7�KK�&�\jD��t��\�j(���(�c&3B�F0�U�	�D�DFTe�RO���ȂJ	�I���ǌ�E6j��7�0b�3N�`'�[�Wh��;,�s�T�`��9�Z����$v�j�d�ֵ~ m��b�?�yt���=���H�U3�?|��|��� Nɫ�3���86�&��/�s.��Q���#����݈b���R�e?�>�	����<�^���;������Yz����q�߾\���e�`'lm��h�t�%�J3�%���7>K2���MD�����7.�e�J�|����[g#w��!`Ճ�[���ѽe��y3+���n?�8q╚��1N�����7�v͒'���<�\�ںD��<'<�1n�E�e���v��Ľ}oz�0:]Ks:��c���_��0��l��T2,եݯ�4gꪤ�)�7��'����ڊ�����4p�ɟǙg����į~�+�*��}%��;�?f�լ	�S���S��e�P2D�8��b�n"���yI�=�>9���*�n=���N1���T�JǞԯ"�����&�V�;�Ԙ�'$>�t��|�ny�0���Y#L��Q��6C��)�GA[w%73�R
�J�K��.�W��^,QM:��l\Lc^�[�'K���/�t�������k�H
�H�38��)@�U�9D��=�R��ظ �@�0D'i��X�ȹ�`�62�*�C}�8^c� �6/T�2�ԛ[&,ʳ� �`Foڷ!,Y���T�@@#�w�G�]�G�@h��"�kn��3���@1�xMJ��N=!���m�SL�fChq�t��lܡdR�6iY�����"!#���%�X&��Uh�K瞅�/:O�̅�=�?��n�����m�.��_�!�t4.o�/��^|e���[/'+1�llX��&�gr��t� ΍��2}�r��'�Nu��+�M�U�q�"� ���d����y���zy�qs�����ݥ&�����g��Ǐ������O�--Ff��w���Wr�y��<���ljW�m��n�v�mbn"����5ע3�C��(y]����<'ժ�p�c�5���j5q�0d��ƕ�]r$��aױ;ᜳO���%���}������XF7��7�n�M�ގg�x~�����2qb� ڶ��"YOP��1��!�J�yÂQ	Ii�C��t��^���*�BYƈ+���ĕ�l�D�e���	�h1��p)U4D���e^iQfh<�k#��<�$��0#.����]���X�j�KWe��7snKE�Lr�iNpI� �(Vv8|o����
hh�m�3Fe��S�-^�dg�\T@6T���-�[RN"0b9����c}Zަ���;�/�nS�+�|8����J�����de��j�La0hL�	P�b�	49��aIB�����3���X�p�i�	���%ޫ���J�bB"Vt��'R�����D~�*�����}㤟�獵���auXN=�,|�ӑ\�BG���%KQ(0b�`)��v�<����ᎿL���q��ӊ��ak�ĩ�^$���i��;��7Ȯ�;ʋ��*W���sԡ����{}�^��a�	Q!��	ąfA4s��;n��0�Q�_5%q����M�7�T�~G�ٜ�?�������~�����gp�v�%�y��G���#�1��(?&����O�̯g�O6�8t�Zj�����'`���XR1��C�����8Nx*�Ke��}���	M1X�_�OM��H30�ީ�t��X��!e1vJsB�"�D��Rİ����ž{�)F���+��A�1*eO���t+[������G�!L��l�Aw" -F�ޝz���OзҮ�i���}�C�v	�<��>���@�{ɓɾl�=���^��J[����MpD�1.	��@�.`�0�����d�S~�q2f�2P�
R�MOV�U`T�8i��J�r�dM��bҾ�d�Ye������\o�IDV��k"�c�#�X��&Y�w�~��J?32�| U ���u��ܩ$��Q�OF0	�����D@���׊���a�Y*⩾��� .��_	,��F�qR +]XL�*�KI�,l�9�>p?y�)����{��X�E�f9�0a�f�B��R��P�h,��L�A[VJ��]�<NF��G� ������L�Iyo��E�) N�?�if�-F�7�)�q��g�?.:��-�#�xU�u$�����/�v��%���j"�5q�{��ضr&���|���XQL&��I��wQ`N1�Z��	 *f��Nƀ�ېWWAl��ǃ�ƌ��9��'}UO,��7l�c/��.���d�<���Ǐ�������o ��H߶YA��^��������@��J�NXz��I��]i����es��-���J��8�-2ػ�/]}Zm�cȃ_�b��� .�8ߺA�t*R��nʈ�ﮔL#��!Q��<�0��#1ᨣ�������
ޯpR�!054�Y�ΖLZ/0|o���#s	�+��a�h�?4I�IHx"�%��}�^@�ퟯ�M�u�>�S�9��Tϔn��=�E#�jպ}�z"DW&���KCBک���n˙n6V��YAw���UU�f��OQvh��4i�,�@R:է�T��.�Zv<��J��j�=���;0�l�X�>b��@5��C�َH�T�O��+ݷ԰V��_�~��Z�%�UOO1=7�']f^+|�t˪g#�7�KS�O��IK�Bh( b�L��6z�)u�+o6���#�E�b��3��l*�]UQ����~�t�89.u}o��?0��#g��/_ptJ@�P ��$��ip�,���y��:s���,�z���&��aZ��]IE�[bw�\�z(F-+�`꽗W��b�-��r*.1-��{?e9�F����{#`�!�cؑ�EU@BI^s��*Ïa�~���7��1�=Hd �J��)=��;��߭� ��Me����{g�����'N��F�f��fqӿ�+�<��,�Dc
��z"F�Uc*����|�ϴ������zH�����nYXj��mw\|�5X�fr�聬j9��Qჿ{�}���"J�=�e℡cǣ-Rrq �<ئ2ɻ6��@L�0�R{2�k�!O��8�����B�V	�%6g���@wT.A�r�*SS�.���i@J���nE�E4,N�)#&"q

�t3
R�������l��m����2���W����P�[�d���d�zvOg��=ݟ��.���
��d������Ԟ+����m�]�Y�R�����8�}�=Y9�eQrQ:��ݦzơ��M&��|:��`7mT�ޫ4C�>�h���_�E&X����P ����L���Oj�L?�0��_�����5�rΞ��}�g�~��|�Q%R5@�>����)�ń4c�-f�i�7
ı���z���9��ĵ���-�X�f�4�9��~�u�.8�s�}�9{���f̘5~*{vsJ���M9d�2=�h1" N����X�{��^˹_���rs`�Nڱ��^�P�*J�i>8�T'�fu�l�O�ߞB[�    IDAT��l� .�eM\� ��g6�����F�za���,G�]&�z; ��d�nW���i�ll���+�=���������4�DnF9Y,�ێ��)3��k�[:M�	�'e/���'���ϭ��:m�i!�����נ�uRk�E�Ss��b&B%�O'�M`�?�����8JЕ�؊�߈ .�P[�������J �1G�	��+���ԩ�\��Q�3xz�ƥ+м�E�G��Ϡ\L��[9U��N��p�.GaZ�D 'J)5
�K���>��!:8��~\�;T6��N��ʰ�?��_�]=`�a���<���Ƭ�*� @U"Bz�̑b�R#�^��/tx�
�oم,[D�9=����Cԣ���A؋��0Ş���;�X%�_�P{K
2ƲW^7ϕ�^�6��
H�J>y�<���n^<��8+�F'�M��Y�_L�(���e����TC�Ʊ�����=�4��(�9�=����hLۻ/�y*.:�L�2�����I����N�����>}�~�n� �Ԫ��Gq�EӚ�p,�Dm!��saKf��q�Dh]������.�G8-F�8R���,ح���f ��6v�<J��r0@��������!x��A����Ryb��0�PK+�z.v{�z�9���k|��A�۟�de�{��/�8���-}��z�ɫf͸���j�8
m�z=fw��[l�J��>�"������Q6u,��s\�{��خhÂ��RZ�P:Sʹ�O�oz�Y��C�c�u�X^����l��r-��G���'�}��C�U��v��填�K�^�C�����Y4qll����U�=�v=e*3�������*���$j��Do�)כk,�~sobMr��ěz +ņ�b,��`@��ކi�����~��s5Qt����0�]�����^��
�4�/`[�ح�����ÙY��G&� N����b�TF''+��lu�k�ެ+�F�I\�wU��I4�1q�>*���+�*@��l�u�6e��'m��N����>_�J�J�˳�(hӠ�sϟ��Р�\�T�F���~���4�~)x�<��t�t�Q��<����@ �#�S���/���a�>?e�����]S�-�����Z�[fB V���kADpޮ��L�5�k3��S��lʉ)��<GF�TS�;��197�eF�泗������IY�����@ɏ�f$��p�)�q��_F.G�o������xe��䕔��Rl��ϻ1���_޼~)&N�񕫮�j[�k��2y-������
��6޾yR�)Y���3c�	�x?�Ax��:���ϠP/�5;>i�^]�� i��NL�?�<�
�:�+ߩ�3q�vحg�y�MI���\����޲l[��ʳb@3P�,tg�n/{/�{��Ti~��O�js���]u�xNV�j:]DT�oʼ��F��EOz]�v�G�ı�,��R1!K�[��A��c睍�!�K�����m�W�F�F��SfH����дG��s�����8���ĆSRǞ8����_�TVD�M��r��S��b� 
P�쩤*T�=�=�<_.�
"�헦|��K������ۦ˹r'.3W¾U아��%be��&Q����IT:嫣�,��cU�YJ%-=u��rRR ��8��V���Q�Vg��L]Fd�xFO��iR����q�A^�X�,׎�Z��l�Ѣ Ųm
+�Q[�V���b�������� $�T��bˈ�P��$��A�wB����~_��J�O����ĝw�k76��*��kC�����Ο�Wc�8���v����ţ�?���d~�����p����=q���^|�ֲ��~�KC��|��Y�hU���2���\�+#)v8U�����^�M����)���x�Ή��5(�=1Y�M�B3qø���+��[o��5�DU�$�8�~��j�^��u(�uF���?إ�ON��8∟\t�E7q�]s'�	��S{⸿���/_?��'�Y�<�Z+ ͫs%�M���Ͽ��I6q��Ο:ډ��U;ɡ���p��nEl椱W��f���l>-Yp��=D����Sw���������q2���J͋#e���f0�o/��KE�2�d�����M�|�)�4�	�G�Z�ı����E�qd���Qv*A��9�>qd,mĩ��;�]�lA��4�@�%>J¥:�m�A�B^��݁�dM)�Kc�:X�
�H��\.�U��)�a��X��$�Ȧ��fI�5U�@nk;�����R��S�C�� AZSP�2R���0���T�� Rc��� ^��L�����ˀNﵶ�P���:�z_�H��:����f��!U��Sm7�ؼ�!Iϭ�IT�^}o�g��V.��q/3�j|;�]���ߺ\Ne���q���/Ug� ��$n��/�^J�[�"胟��ؿ� �����{��i�=)`B���1D�S��c�ԵCn�i���ϓ���|��_;��O`d��H��'��u��-�i�fڿ!G���	���Lf�S�Ο|=}_B��Y��!ҥ����:�	�w�����]�Z�]U�{`��^o����89��,���g�C����b��x�ݕ���~�W_}�u#F�PO�Ѳ�A�o���|��i?�I��e>�r�'U�U��rO�O�Pܱ?�
�����?_��Q(%J�G�T�F̜�20b[̙Y���8�0b�6��Y�����lt�=�e����[��ނ��W��(c�hR˧K�&��!����T�f"b����	�3�Q�A�<�
�$0%U*5��7J�s�I�#ؽ��{�L>�@���>���ҋ�^�I^1U�o�%PQ��t�7�릍�U��ڮz�V��::L�3��1=����s��A��K���v��7�����0�)�� �<f
�V�}���l�������-U^V��
0:����'��Ӝ���+�s�C�M�nv�K�H�^�F"�e�� \�L���P�hW���ɾ���I��yJ5�}��`!�Y���6�6��ؘ���q�Tx��U�*��	������B�'�G�����[ŀxP�>8��p�g.Du6���ďy^xevG ;��8W�XJu��:�T0ʰ�uÆx�_~u��_�����͝���~�����`��l]??*����ʱ���5m��}�~�w�X�@˲�",IU������S�U�����/Gy�]�]wݿ6�J��j�� �w?���/͚�CF�����T��\�0L�7��{�[��.�}�2��)ʠ߾���܂(r��o_��Jn 6��K��.2qI�v�%ղJuW��1qb��Я����ټ<�m��ɉ�;Y�1cNSNF>�U����/y�:�L�oڌG/�8G@!��������'c�݄�J<�*���u8-O�U���N)�u|):�8U�T�45��J�e�ِiT��}yw&F�:*0һ��oe�������GEN�E���v�O���r��WL�
 u�Sǣ���ҳf��;4���vb$TT���P@�C
�a���j�E��W�-_d<:�(����,������W�\.��Y�<���O�
z�%L�ݎ�<y3�'�2�i๘k��j^L�b<V��c;Dz\e�V�ӳPa���Q�X}d� ���9T�!�^���d<��(>q_��e�/�;�p�R��c����5�9�`�U9�JJv�����{~�E˗�*��F&N���	��A��(hٲ~s<�Ͽ��ߜ�ہ�w��$1�̙��;wn�9s��7oޘ�k���y�  �M�l@ϧ�����޻-�
�;�~��7~$�S���~�3�w���I9����H. �c�v�5ڱ�wz���V-��?��;��8i'�r�7]6���ҺA���%7�.�cv�Qo��4��2prH��������_p�g.Fc�8Up`�L`6�nC3~~�]x���`X.Z�ې�g� �}�{�hg�$@�RN�[��S����F���a塎�C}�^�jNF�$�Ƶ��ޡUƬdش'��W��A8�@���L$H��d\QE?*��%{B���f�j�%�k1�l/N�����R��i����ۂ1eE�X@1���W��xd�x�I2�n�O{�ԑ��P�J�@���\�X�\����� L�VZ*���%�롄&��_=�����tҘ���Ʉ̂�o^I�S�����s�e��X1O��)�&�
�Geu
(�x#���>q��0"[��}�DF��#�렒�(��;��T� {I}��R=P�k4�2҇�TV���凐�a�$	"�E�u���p���Tęm����R��*�:�B>��8&Q�� ��Z���{?��H�Oi��G	�:���� �W^10LΡ�QX�~g�Q�Ŏ���>A���6`�?��k_����r}3gά�={v�Y�f��7o�	A1Ms�eY�I��Q�i��!Ho_�����l�<�"~��iZZ��$�a�0\}ꩧ�x��w?�A��{��N��~����楿�����E�eE���m���W4����!�����kw��q���o|'��ig�#��P�騒��8u��w�/��q��/�i�/=�tx=�ck�����/c�aC�ګ�`��O˵|���c��!x��9�凷�����E����#gIx��R�edA\�׆S���RN-�8u<��a�t�Rdy<*�+���;:��?j�M5,��� |�6I�e�!=y�m�{���4HTO
����H��$9&#���E�a}z�$Z~�Г�Re*�[Q��&\2y���Լ��<�b�
l�\Y2S��gУ-A.P��c�A�]Q�v'���wj�(B��<o�p����R�'uf$��9LY����%[ـd�����Zٖ���>�����22t1���{9� V �6#bm���q�C?�����^/�D��
Ta���z|Ӌ.�
:���gO1��i`M����p���-�I�.�Hrj��3n쥸����md��k�b�I~����Z��S񧉓P�T9W��e�ɞ�4߰q&O�|�	7_�=�aw��w��{�ܹ�W�X�@� be�GY��\H^Δ�������1�h4R3�r������@�J��[�ap��NA���;��o��&u��͖����������SߏKm��Fl۶�A`v��2�I��DTJ禞D�� ��i(��0���`�+�PѤ�`�Ru��@Q�m���+�Ի�}[5���?{������N���x+ǅ�)�~�56�ĈY7Bl�����-���5�$u�{9��	�ܫ���a�����Cd���i1N��˃���1 ΐ�]�W�mK���%]����'?�	�/]&c��Ѐ��[X�����4{� ���"�iz	 �ĕ�� �:ʂ���mAܶ��2A�W�Ti�ə� ZH2�J4pc��@@�Lw���K̅9p"2 	�QO���U�b�b˃�D�H�M�0h�+ !Mb(���ϯj�'H"�t�HϦ�2�U��d�kU,������*���+�[Pjv���r��D$O%��h��œ�BE��U·�EH �Ne��S���Q���+Z�O�]��xd��8t�WeV����rT�}[F��r��:w@Q��b圦%SI�H/�N�z��Hߨ�z��(۷l�m�+ NxU��0n�e���ߑ�� �3{�/]�?�e2��1-�'}@��M�1i��;&L�o�{.�?�g��Nq'Nt��{f+�����Z�/
��J���1��`�5b$	�բ�4"yP����2�8��2�Sy�n Ӳ3��G3�]�cc���ښ-������\��r��ifad[J�[
�Ǒ�Э'����^7+�����v*/+���<����G�+�#�fY���?L�Z�c>�$@l8���65���l��7�4a'!FF��P��I���x4A�E ��_����,��g��Ŀ�Izh$�����+.���8�!������W���յU(A��~ N�gEy��˫Tv�U+J`�,[;Ғj�U�D)3E}���rK��K���	A���b��b����V�yg�D���Yj��0"�1�����<:��a��g1��=�����Y6~3	�ĥ
P-P�)�o'b�2M���J�Ņ1W\?Y;�#��*+��Y
��u��t}d����G�a� �)����s}l��%��1ZqF
�d4d�JS��
�qP)���S%(�����Rʿ)��u#�8� b�t6P�~J�.ה����[���{�+�b��*����m�Q#1r����K68��'U�=z���M[���s�r�Z�J��SN-D*�-V6{�ʁb�&����7����v�+��� ��8h�c�7��~�>��O.��3��J�v��,a)b���
$��|���c�u&NGҨ�K�����k�+��;>q���4������u��6z64�_�"F~~�Q���{T��rD>B'��%�ʩU,��=q���Ľ�q�*o���/}e)��*�)0���էT��#.Ʌ���_�$�Hu��<(�v	�V�T.R&M�;���ؑ%}d1�K�{U�M����s�F@_;�yM�o��O]����O�S�� �4�f�j�N�i����U�1 )��]�E�bg��V��U|e!������\��0�T�,�+(*�>��a�0�G��@U`M��)捋����LVud �~������rTuKQ�U�u }e�R�!U��T�Uz_KW@����RU��(�\Q��E�*N�u�[pW>�'\�v�'�SS�{�?����_'���{�t��=�v� �-������򪫮9/��K��H�YJ���j{�����.���8![*z�䈴�2���K/�|�c�:��<�����r8x�A����k׷�?����&�������^�|� �ҚG��J���+�:
��Y�K{�ҙ]#���l"����u��J��e�����zה��R��^J����T%X��� �b OT��������FEIR-`���&	�����H
A�����8Z\��u�"=��=��\��"p�lI-`8f*�^5�q�t+`��
,�Jy������	%�G�b�Z5�$"�Oٗ'L���S�Ųi&N�l��%�b�`�=p�JA�\��q��B�y�rZH��J\~S�o�O����
��8m*J=�����;�:Lb�ݲm}m�u2uՇ���S��y߸i}8q��}�k�o޾3���=u�Aܞz�v�~/\�p��z���Sxcc/\F�]��D(�����! qRO{��i�G1qI���נ����)cF��Ԋ��PU�G�>�ز��3O��O~~;�Z<TU�K�3c6�'	2�m�`�h1rJ��R�5&�sSY�ZfLW��ߛ��$q���֔Q���/jR.���K�&.�㓌�X��,�*��ʉ
pH��ʉ�͒��W�aI�q��#2�JS1`�0���+k��f/�%�A R�*�JO��)vP��	���(,m���5�%
WQ���mҫz�~)�ƅ N"��rR"�:|�R�� -��!�xP`���t&��i�k�0������D���x� 3�2��Ɛ��q;�mUcePO��:?�L+0[5ft��ȧR#e�
f�����Q�A�i!�P��ǩ��L�����K���Q��R�
�K["�T&�_&��M냉'�򵯍��v����#������v�����7eʣ�7v���Ea7�lyx�#�m/�e�> �	��KTWg��Qd�3���?g�u��o?�jh�۴e3^}�U<���X�z=3#|
K9,�~� N)P�5�G�?��i�@=_��Fp)&�=���#�>�\�� +}bL��N�K�05C�{ܴE����N�VʎC�V	���,��V	��J���?#
V.>�R��O�����6ո�X@� ��U0.�g%��7�TaU��hm���Ob�(�RecզJ�ơYeUR���DQ�$U�J/`$1^�����u�2�>G\�l�B	AW=}�u�j�P}�ȩ�0s����K�cU��Z����ە�u.�����S�Ob%���e3�uMX_�    IDATs�Aʶ�X=O��C��r�x�U���i�T�6l\L�<�&L��[;jn�^Ϟ1� n�8O;m/.[8|�C�=�WK&���DfWj�9E�ѥ�[O�Eɇ��#�t2c�'<2>�7c#�=������~d�X�t	V�\Ic9�oP
�L�Z��^P�A����ĩ�t��P���ypr�q�K�l؈O"��S'bDq�T���|"07�X@��]%�;���Y��\�YD{�g�Q�C4�<��*d��q2��
����vK�0�N�B{	��zxq�����El���� y'#���\x��fzP���U�p�=G��f��M�lӁ���X�-����c���FB��؂k��"߈Qby�*�5m8���$�a��B�u-X~A|0%3W<�\��K�f�Hl�&��Vq� F[�����f��ᢑ-���39쳤�WgM[<_<�9;ۧ��7�ױ�kٵ��az��
�NB@;g���E���C�vF�_��X$eX�K���,���Tt�q۩�L�#S�����pSQV�o�{��,�N�<������ݝ6Yt�x��n�[��n�-Zt�����|�U�)���h����8���&�o~]���أܞ�8����I���	���M�ͤ�X���l���з��wǶ��k�a�����7W�B1�u檲(���
�e�;�8U�SyŜ�Mq��`8����0B&SE�a��E�#CnG�
L$N-��4P���V\~>����0��H
��� g��cD_���*����Q�������	-\8�V�[d��a\Pi��
Eaʦ�	�r��.R$�6���dVq�?��իQ�|���V؎��_D.�E)��1{ӴPc*�k�b#A�*�R� ̘k�ȘJ��b�!��*�����fyهmD�0�	;�
��x4O����xTӅ�kN�CF�b�v6�@�$HU�1m�12.��!ǅ ZCs����"A0��4�)�%2Mv΁/}�*�0��	�f�hn�"����*�����P��d2��)؈��R�UiUXXծ����Q�W*�ٖQ/۩�Yj�J�c���U��I�&}c���c��k��G����gh'�A�����7��*A��cf�
�%:����x�}T;y7����I�9'����!�@��qL���q�QG��~��=��5�P|���{�F�,Y���{?�MT@�;�͒rj&ީ���qSz��JM�wdv�X�}""�d��%�Ā��c�U�3F6IPl+©�����ճ��P̄(2�#��ұ��.��[�a,�=HJf �U�������c�)m[ȆY���ȹ@\���`#�0���� Z��@��v��sa#j)�6GIf;נm��ʦ&�D� ״��_���P����
+���*��+�0�Y�2�����\�.Ԓ�)�����z@��e�Z�\��q���"�lfU-�v�ࢊ��oU�~'_����i�0�6T�L�Q�C9A� YZӔJ�MC��Ű��e�1-��)�,@����hv��M����V�Y !B�:>"�G�l����}��*��,�$=�d m��~G2�R|E�{�z��[v�S(S���A\�K=�iS��?4 .�<y������`��F�'�����oO<��}�v�\�d���<x׸�W��QN%# �A��9[9��ߩ�h����NP<�Ī�JWw���>�{��s��'?�q��V�D��������QWS��{={��I'��^�����,_�Q�J�?�v��HgW���1	X�c��T+�z�����!bx>6,Y�⪥ȑ��M��{���0�9#D{Ƈݳ/��$�ڞD3�[ZT�_������r�>�q���>�:��߀������Ep�f��˱�-��A���,��z�7�{ �� ?B��	k�BӊŨ�6!g�Pi���-Rwd�Ȁ��yb0Vߓ\���X&Z�C;ց����B��^�j�'Ah0:,R�I<N6���\\fqF�&>���B�������c3�]߄z�'h�K[��F�a���-�"غ~܎�k��aG"Oe��X;w.y.�%ӂa;�XCD%�|p�6��Z��8�c��������L��}đ	�Ȫ��$���0�V�f`���J@^�gy<��R,m6E����A\*P!���@����&�z&N0^�h���U�{�����#��i���?�-n��;�@7����z����ŋ��:m�/ǎ�b�b�Tແ8� �+�;;vD��E����T�I�CC�:�`���?����7^�������G~w�}7jjj$����[o�)f<�<"*!m'���S�~� .���(*�He�H�Ӑ�*��3T�h@�G����S�r��|�.��X8����ig`��c˳���}4g|uϾp��\-�ڪ��V�ĦO`��7`�#/c!���p�
/䀪:�eZ����/=�|1@5!���hf������c`z �#���Œ�Z"x/���'�۶	~d"�V!�T	�"��,A\ ǾI)�/��ZUH�K�gG\펅}O>��|�SƲIO���bc��jd;��BS�u(�S1��O�ҋF3�-Q�u��a��ҭ?Ef�*��eO���EԌ�~���%�M��5��"Q[~]5�t0x/`�"����C?�7Жƞe#��B.t��]�[Q��`Y>�c����O�p#�*���<����,,�!���`�$�͋�ȸՈ=a��lƁ�� B&,Q���+��Lemղ���0q�io����o�&s�sO�4�	n����C�{���q{�9��,Z�h��S�|���Fj�X6���ĉû,j���AS��f����4�
$���������~�����Ҵ	?������{�[~���~Z��O�344�į��?�?�1�+B6��Uۉ��R�-l�n�*�^�KX�U��B���{�>p�x��9��f0x���k��ɓ��Ԋc/� 8�d,�6-O�BuT�V��>'�F��.E�ҵx�W��e�w�a�9l�`����0�oDM��x�ɰ<X��g��`�Vę�2�#漀����u+2x��#l�N<s"�|	��6�[���Ő}�Gè〶,���&("�sh�}���	K�qP(�zO�� ��U-��*;As�~m55
}�]�uNǚIO������`���h���8�(����"�|5򡅰��99k��~����`��|=WoF�I؊$�`��A��c��_�Jއ�3g I	���aW^���\�g���iނ������!�B��,������8��������|������7��4�>"ۅҋ�E�� ��E��[��h�b)�6�r[�"k$2~�"q�2qi�ٶ�m=��w�.���>T.����q�m��ߵ��@7�����N�C��M{x�]��]q�0q��`�4�S,�,�����@L[�{1��V�2Y����?7~�Z<;�E��$���	��c��~���_ㅿ�(Lܵ�^���������8�:1;5r)�n�����>58=�5�86��R�BYw�G���9�"���%@.S_�}��0�h̘�(��8�cg��IAXp�?�xV=���?��R-��a'�A��K���\,y�>��k{��s��=͏>�����}�G�/_	,]�~���dC4y����a��Co-`��ŨA��k�ݶ�d;p8�~�_��f�l:�%��Ȱ,����?HR������
�W/�y(�:�; X�+_~	��G��	��ꇽ�b�
m����� ��[�~K,�Y_�Q���`�2lx`&j(��m~+��%�l*�9�0��1�?h?u��_��/�������pҵ�
���m��Y�ua1Zd,x5�0���P}�8 ���_��&a���8�̳��� ;����_��V����`k�:�u�p��@�^�Vn��^�9���/�z�t��a�O��'вf2{��~�s�H�ß����������h�m��ы.�xs�$�֭G�D��h�#����S��u��#@�.��}Qe�mAݶI3z��=��/{�:5�4i�W����^�{��Aܞw�v�����!?��]��]~�?q>[�o�����a,�QJ�JD���[��O��㺫E����.��|�c���"����*��؂_�}�=�$��E� .fS��ߺҋ��V>	�3���*�+�NʗEy�b_>��3R�-��lA�ꪰ�Y?����mƨ��#�GAu&�CN;8u�=�8�z��� �`�'�9�3h}����{d
-ؚ��p ������x��?�I'��2+�z��|�a��6�U��b����x�',�Ve�R]�����K.��̳xy�T�moFM������ђɣ�ıt�����1�=�T��
%�ڋ(a�Ca���ػ�����}a[ѣ(FX��(�1|�gS�9��g�&� �
D�v�~������]����x�������f�
���_�aC��-?@�굨��0P@�c�Ի��sp�� ��͛�h�t�;<��K�6lz��������T��}�I�>���g�Ęo���̝�&N��`� ��\�+�k�Z7a�� =�����k�����Wa�����l-��_��P��ȅ1P("KA	�Q�[O�*�b;��ߛSW@�2;V~���Z�/�dv������q���u���n�{��]�
�=r׸�W(�$��8��;��w�n�����8�e���CP!$�^�lg�q���yٶ�&�F�c|���wK���;��c3���Az�H����T�E������>�8=��g�Y� �ta	��-�\`�'	T��(5�%	�e3)@��H�A�0Qʹ�z�a�9�c��!P��6`�cb��^����?up�qX7�Yl�w*�"|7D���E���������Q�҂ �bSM-���G@�3���v����ñp��h�q�<i�c�e�^D�*�D[J8q��C�>�s�	h8�t4O}o=��[7�����KU��������>��K���!��쓁b�M�& ����=��ş��ͫ0d����+����د�¨#�B�O]�7�xK����9�	'��ŗ����о�N=}>v0�5̜���8�3`}6=�"f?�N��K�C����6lFC��\\B����m2#?y!P�mV�싅S��y�zy�)�#�~>���u'��^B�����WP�7��glY��#���L��{'�*���;�c ����p�G�=�,l�=�=���Z},r���?�Ͻ�w���o����n��7��n߂<K���HDy#�/��L�`E��ĤW��m���u[���q�5Vf�vT*��N8�1�|���ح��7n܈ɓ'~�[��~���{�A܇�<n�Q�_�t�G�r׸�ǝ� n���A~p�@E4�mkkC�u��֖���E�t8�8骧w�<�EK�|U^�$�n&���0��<��$+ ���U��F�c�vı�� �P&��L*�ݷ�&�	 ��� '(�07� l�Á�+���^�Wh����:�{�ϱy�2�|�ǁ�'`��Oa�Sѓ�m�O8֧.ņ�^������V��Uc�e��_��Z��}'�|0�H�y�l�9���֢�Ҕ7��H�@ M~�l��G��O<U'�F��k�>�~�Q�KE1�-lę����-sc�A���u1���\��#�Ɵ��֖���%@d��[�m5j�������g��q�	���x,=2��}:��O��3���ð�?�E`� ������\9���}/���-xm��8r�I���x���v�ZT�4�&	іs�r�p���@K��#�9k֬C��0|V=�����u��x�&O¨�G!{�8ly����d���=p�/��~�s4mY�s���ꃩ7܀��&���R��?�6�>س�J����a�9g s���g����]�|m��?���5+PeyȻ���i���a.���3/v��#�f�Ʈq"l�������┙w�C�ĥ~�w��m���q����=���8��R����Bd�U,T��Vnj�,�o�����'qmL�4Λ⤟��"(��4W��ĉ���<r'�HT��y
B�:(dDuq�9�����#31qʙ'��i��4o.���T�8�TXg���<��i3Pz�l�`��ǡ����ױ��i���(�6�~z]�y����u�O1���/C�����5��r�!�[�6T�נ�y+�,�%X��Bl��A���\,|/L����>I�R؊�)=P
�A�އ�ƫ�������LAc��
8�s������J� c��X�+���I3�����X�gn�_s���\r)�Okg<�cN9	8�l��w"6Ϝ)��C��	hh��w�M˗��d���C/�,�Vļ��@��G�?���ȵ���^!�">C��Zz<;s&�:�l�}zI���s����1��+P�=���-����?3k�{�(��|�/�$p��x���a��U8�7�FL��F���1�ˀL^��$�-_	�T@�q�c��O��S�=���@��'^����o[32I����D��V qN�&.���C�S_�l�EL\�:5�2j�syU��ʩ)�K���o ?L��Ǐ����tB���>� ���k�K�,�롇��9vܸ�>�L{�$~��D�%^p��,{��L�!�d󎓧����$!�Q��d��GMSK��S�8)E1 ��Foqd��X�8Ɛ���7m���^������3ga��8x��=� lz����S8��O '��53f�y�_Q���ۂ��>5�]���'g�*��u�. j��X��Sh�;���7��
��NƖ�����쁁#D��,��r^(���ɢ���o��b�W=6��"6��2�֎���G�^���C�[��/����1�+_��b��G�U�ާ��u2л�<A��d��5�x�緣�SDܫ�~뿀���[��G���bʹiX7�	v����d�_Pz�x���>�/pN8�����_g�y�!G��3�E��l�0m*��̅RN}����[P](�L|�eld�AW\<�{�Q�:�t�:�h�G#�Eoa���D.���7�'�z=����1�o_��s@S��~7oE~�`=�l�.�L�#V�]�����Gn��9�������YX��_�&��9	��#~b��ʫ}�W�����5נo@�� )-a`ñ�h�lW]N%�����mA�<�t|C;3tۂ4�6m3�a q�&M�ڄ	7���5�t����n��Gx7_�[o�5��)��7n��E�"�T�(W9���T�� 9)��2Lz>�zI�ư$Ղ .�d$���t�/�,�>ÝQN-�8�S�ډ���lM0O�?��f��B�wO<�\��Sn܄BSj�"��wލ��&y�E�c��K�[�h�:��3=F����n��p9�hT^q���{'��bs{=�>��;�=`�b�e�7�PLg<�L[	Ái���Z�GÅg��2^��֯�I;��{��^��7�t�Ds��� -RV-�ƍ��k�A@}5ڟ��y/�F.S��.�hjë��%2��@�F���G�-�s?�'u,���bՃ`��'1��3�����B����Z�p����~
��,�/I���<��>��o����`ľ����ת�y�q^Cz���3�A��x������a�������ڇ�J����|���+_����a�>ΨC�yK�o�w��@}�����X]؀Ӿ���3'|٠���{]t���mY8��y����=l��d�X����M �b�~��V���$����ܘe{���k���1�]�Z�v%�a[e�Tصmj��NtT��Im���M�4�[&����|��޽<� n螶�ŋ�2m��Ǝ;�'�    IDAT���$��b����Z,v���R��<Û?�:�e�(�g09`�2����Nqj_��. �����AB�d��{}4�Q�5u���a}ly�Y4-\��1옣a�>��	�֭��Y�ô�4�4���d�D�X=w��,Da�2�W�(&�k����t�)C¬Q^|N���ƿ>�h�Z8^����_�0�5[�欍ܨ������wo��d�as�y+�����X��Tk{⠳N���G���/ �Ԇ��z�{�i�-����HZ�����]}ZV���ɏ������1k^xk^��#�<>�^�����blr]�u�H4�?гN�A������xk��N�CO�9L��x-L�LN��B�#C�a���ٗ�j�R8=�0��c�>0逸�[�HF\6N��������>�8���8��Fk�7�c݌`����*�K/��x���Sl��ǌF�Q#t�ņ,{n��iÒ�}�d������N�Q\���}�fVŅ9��u1��i��#��^m�=����vcه�Ly"�//o��R����&����9ݟ�sG����n��9A�CS����q���Qq��I�V��##G`�ٸ�.U=��ro���S�"�"8L�]����ԭӷ�K�T�&K��C��J�I!M�5g��ˀ�3����͈I���^��X���چzlZ���6pz.1ҩ�Iu=|�km�5m�mfP�cox4�C��[[`�����.�~�\��m~���j���W� Œ���lZ��q(�Pa�#���IL��Cs�C�ς᪍}z�(��7����n�	
�:.��G�8���0��[�`ˊU�Z��,4��M�.o�<
=D��\'F�U���i�$M-�٣Q����&���h�c����5�ٷ"�@{K-M[ �+
Q[�C��
[6l��%�r2O����-�6I*B�Z���ĩBӺ5hK���?Dz�M�el����D��}��l*�b��5ȷQ��h�������vs&U�T�����9���\D��h�Ç�>}�:�K��_���Y����J�� �E��}��%��+�n���J;�2a�!a�n�0��v��н�=f�A�s�vΎ~�A\¨釣�N�ų��y��ΉPH�w~�) ~I�8�]e�;���v�=E�b�@�n��b��#��:��n��J��2�c(9���Qǐy&��`H���͡�}�Q�\���TjG�e�B;�rY)����$!�l��l��"�+�A�������6	f�|o����-���f�����_�-=�A���|�W@��7*w\π�R"��]�yJI�ua[������h��X��N��A�ж��7 �'����C�fC%!ۀk�KWt9W����!rD�ɒWFTyv,���J�k��w�(�(AƭEk[ׂm%0�2�!��Ҧ�Q�c��2��Gbǒ�J����Dֶ`�����c�k��vs�=X����3.���a�R�� pc#����k�k�0�,�8����&��\˖8mp�l�0=��JD���i��GpaKY�L\hR�$���tW�L]a�TRIgP�>N��]*�����!q�N�p��]9ݟ��F���y�l��1{��2���*'��
6ͼu��ӲKy�;��/�r���V��uS Td0l]��uq�#]qz���$�@�0���#S�E$�B��N��^�V�r� �x)�jV�@����(�a��/�#�ʶ�C�D8q�2AF���j�#���y��v�FH�+�yq�,���X�s�-��(���\�7�ӄ���s{d ̈́L�	ߴ&\�S
R�~�x�X���W")*�R:=���t��c�Y�Oj��t�RE���9��{!�u�{]�X:s��}<�X\�Z���E%$�}M��"G�8��Vۉ�$��S��,wl�7�-[��}�&
.ˡʊ�c���^Eڽ0���^Σ2�uBW�DǺ��0�O嵤�{���8�=��+�?%�.�9Ð|(�o)�h,��$Ɲ�����k�|2a�וd��MAm�� �W^10LJ�<���!_�t�;�F�.+�-�R	[�n������o��|�����3� n�9�dO�N%�����u�i�����m��c@�Kj� s=A����z��Z1x�
��� �&{���(0C����*%���4�������A\l˄O�Y����}&J̕5�`!�]���b�h#�,�[q��E��D��eI"��Rr,��PgÊ,81�A����|���I'ce�!�U�昄t!&�J�FV�O ��	|���/L����QA4�Mb�b��c&��1E��
'�L.�~�@W��IMi	���
ʀ IV=(�:�1�Cz��c�^�bd		���Ehm.Ac�✘�(�hӦ�4'�$��X�}��2��MG9vkׂ82��
�A��EXf�@����4�N6\N�IƝ<|8Q N�[�SW�ZvW�	�`�%����g7�t×w�Dҽ�]6� n����7�\6��G����N}7���;�k���^!24������i�c��lN���\���{zPQ
��|��dN`Ap�&p~� �#Ҡ
5'dw�3B6�,IM)#�QrB��yJ�k�+L��>�}hEj=*�W�R�T�L�b���yT���l�,Ya���)cc���%�,�E)
��B�g�Jr&[0MB8��c'`���cx6��7��8��#�J��\��f
����+��Tt���$@
S�(^7e�У��/6�r��������ܹܫ����D&�7�I�SF���r�C�}�K<^7AO��	z�)�+����m�CSZl����E��ݡ~U�GP���eK����4��iO�j�]���C�є|�:�+�&f%���P�JjM嵻�8Ƕ�x֯_�{�|��	㿸{�,;~/�D�tq�|��k,#?�z�)������r�뺆m��ϲ,c�ƍ��%dY�i2{���q������#��(4h�r}��n���r�/^��)�o��&6�8����q��j�S�~c�ԇt��γL{�R�&^�dJ�(0i��R	��n����2c���  �P1L��S,(����ʩd��Gbz�T��3�y�<;g$t'SehAI�:����qߥ�Kƅ�� C;�o$�XɈ�?�2@f�%��R���]d�8a-=l�^E�Щ-�+A�g+�Xn��u�;Q�⒭@S&�K(�kn�L �4�����w)��	%r�1#���23?� �J�};��S@����S�kq<�?�*
�H���PL���P� R�A�r˯����ݮe�ہ��(����ʘ	2p�b	�t�f��}�������q�j0�A�0si����ı����n�:�w߽����&|ნ?vֶ-ZT�t��>�<�̠-[�����Ǳc��EQlF캮��$�a��-��$O��r�&�S����ʿ��|B�?y�M�$N�ĳ,k�!��o�q��:ޮ���ue�>�}뭷�{hʴ;ƍw�GQ��-xz�����{ �R��� NB�;�!50�[��J�^y�-O�z��_<�T҃�q餟����n�%�N�CE3X�,�K@6�Q��	�EvO��q�21��b{�B투��v�8�0� �Sf�~1Ó�L�.z�4��eG�'y)���i��bf�Q�m*�@���,7<�����eb��\`	[�I���M�iY.V� r��49�̖� A��E��]� �):"0�M�c*�)�l�8�5�Tjd�ۨ��XW,�*s�,���r��+�}SW��F���:ʹɫ��^t�}�ߙ�'���Q7���b
����"�SS������M�GbB<��A\��=��#��d2شi���?����n��+�cW~v޼y{=��{-X�����׏ܼy��Q���G9˲��u�f�~杳�I�4u�Q���2d���-� n7:�bW��~��qcO�q�sv!�KK`
̨FsU2e���O�y_�/��d�J9]"c���8�-#U���@��@�a�gN�{RVe���T�H�	A��U%A�<(,�^I��[Ȅ��^�a��K�����r�쥣h"$�'�C�����\+�iyW�K5N�"\(I��3�қ'�'2�)A�)��+גC�28��d�ܐ�#�T�_���0�9ُ,e��Dp@@@�M�8N�S��P��qqS�M̦�3i�ׂ�^)]�M�,����X�r<d�ɤ��iP�ǦK�����5]���AaY˽�j��uVVv�:&N�/'#��(��f$�7�|Q(s\;�����^.T3s�)�!C,f܊	��=�E�AܤI�~���O�����v�g^~�e'������f�I{{�Pg����+�/�����_��͛7����^ EQT+�9��I��A�\�b��N��w4Z�r�a�M���x�СC�w��w̚�A܎�=v-RN�6��qcǍ�qo?�:��O�(w=�ӽB��M@Z��J����zEʊbI��Z�V��b=A����F�B5��h���i�aG�q9��C�(��R&��
m.�.�ٓ���s�,��Z�4<�eM�a	�~�i�D�=�(��U�d�B]O���^1��P�!�3��rf(&�RD#��yV>��	S�HU1���h��ghy���*aEv��>ra#��9�CG3@�Q���\Kd&9��b�Fy����^:�i�J�2^d	�W�by|i���2�ݣ�X	3�`A4*2Y��Dً����V%c2w�@�,{�������Z��k��F����'�fG�
U���m��}��ŠAq���!����֮]�o.�򕫔���A'��@0-��_h/�����đm$��8q�wǏ����d4k֬��r�����9�SǱ�$IE˘v.��y�����8U<�7����� tͶIy���Tes�]G&n�1�u��o��q�ܗ�#GN���>w���&����v���+ve���{�?��?s�U�Ŕv��<Tw�"1���;�/�w�M�Ǡ�����ꌒ'k���%J���O���������)��L�NjP�j
DUZ��=f&YeY`�'˰�D!�� �'N��v��*�����'b[�
�U��N!溇NEwq�	6���J����� ��b����t��L��֥O{�L�+
����+V��Ԁ,����x��^����"�+Ɉ9
��8� N�=���>�JU@���k|+Ab���,=&ҋ��aOY@�9�K
T��KQ����sO��\�CG�G�|�3dO�T�	Ɣ A��<���Ci�B�3R=w{�W������)�) M�]Z�p!$p �*m�Z���'FGu�bX�E�l��,�W���kL�p�*l�sf��Ƽ��S�E����4#��_um���g;�0@6gcԡ#q��g�#�@m�*������۵�[0c�<:c��X���n�J��Nf�3"}U���}����+����.����a����;s���\*��(eGt����4;5��&~���,}��Xl���������[��d�:X�S��/[�l�o~��f�ّAXZPB�20Sqt�"��g�Ә�fߤ�1��ѯ�l&����r�!���/]�;
�A\�<�Q��������³w�x��S�l9�J:��|�%���L���)��j"W f�X��qRP7mu�t<�a8NF�M���`9�f��
"�cK˚LL ["�A��	ĵ�f�]6��������|iR�͔0A1O21J������ c��C+G��bX������ ���ӛ��:�����\YaDxCg���80X*
"�dr�e9��=�`V�	2��6YEy�P0��U#LJ0h��Dp���|ئ�Z?�+"��4��l	�(F�f`d�bQ$�#4LZ�d�g��*�7!�:hlNQ�!�ZV9ɴ(����PhiFUM�C)�Q���UP�D�h�
�
���$�X��Wԯ��)����\w��TTW��Tg(��I�*�׉�ʖ3�֗�~XI3�{�Ρ������\D��=d���ԩ�^����H� �.y	rn~ɃPW�G���ʢ_�^����řg���|F�%�7��H5
b���-�[q�}bƌYX�d92�js�^Ő:R)'�(��J�|��C�8|����]�'��0D���o}sޢ�������.�ǟigN��d��4�{%JQ@�^;*6T���W��Xl��^J��J�AD:	��J��zΙ3��y�����&!ɲ���L>�9ٳsf�3������<k�n!��u䈣4-$�̈��]�-"�+�E�O\W�[����LƟ�[��NQ!4D+�����5M2nܸ�m���[1`{�����^�J�y]�p�Mg�u��M��R�hI@\���m�M1��FS)��z��ᆺ�;l{
�&�:B<ia�_=]�?�T�������,��/)�O�J�?#������u {��5��3�b �I�9eLs/o�>��֦�ϸ�['�,7��c>��,�)ތ�ū���z�(���C⨪O������:�p�u�Q��O��$s"�Z�q�:q��v� ������bS#��䢇?�Ef�L~&�TM�T����ցR[��]��\�N�5�fQ6�C���<�b	��	h��Än�rNP��i>���\��MG�PB����z:{h%�M�d3C��bs�7^'rV��):���2����m�ğ���W�B���JTu哰�g�SB�N�;:T�:�u�
�Z6���VA��tx(b�ՙ1l�H���47B�Bq^�h���������A���r�CH�Z�㤊e�>?��o��Jf)�dZX���^tB�|�u�ySb�Ag�0��ti]üY3���|�;W�Vp�|/D>_@:�E:���2����u�?��߱l��x���(]X��@��JO��!�-���9����s?�@�ÈO����o9�����֮]K�Q�G�:���:&N�(���l<.�7�^�q��Uw8��۳�*�?q��G���w�Ɔú��n9f���ߠ��>ɳL�/�f��)ͧɠ^�t�p�e�'3N��i����;��{���������(V^�k���)m��|��	m�^uՑf
Z�
r\�#%vq�Р�}QN雓�;'��̱�g&.5Xr�:�n�cGb��P��;$ �݀��S{�n17�f��e��7���V${�Di�K�X��P�P�PL���b��Y{�q��ɀ^������V>�f��	�~7�Eo*2@G+ܗ^Ʈ?��歨�d�p��5�����9	�a(����!��Ӏ���\��<���9N<	�9I]��6a��B��0�ԑw����'�渷�v��GA�[��q�QǠ��MMX��_��6�_*3���y�6���ǟ@j�&T�.�B;�29�%a�.Wz�B�G8�
��30��Ӏ�[�����<X%)χ͉]�4�ݪ���d)o���#����B��k�8�@Q<J����
��<�ϰp�\|��Ǜ���'�r��-�76cͺuhilESS2���*Q;b8�L���
vQ�ы��?>�(n��6�ߴ	�I�#k��N��k׮�b��c�:ujX��o��+w��?z��<�����g���	���3v�����޼���Z��Y7ƲR���iY�>���C]��D��p��:�bK�޾*n����Μ�'�)xG����t|�f�W�i�x[3�[�ţr��QW��.���IT\) ���f��U%߇n��DPc#�.G^�Rz�'.�N-��ѕ��I�Hl$Y5(+i�0L4�r�&c�g �#Q�u;4�B��@k���_C�-,��W�^iX�C�T�,��?�'��|V��!�2UBt]X)���U��g������?ؾ;n��[v`f�B���Ђ"�L<��-�#��v6� U3fa��?B�v.�����7Cd'M��O������\�!ë1��W �t�[�\eP3��;�����_�f\��@�RB=̣�Ԡ�����{/�}�<� Lׄ�Y�k��L���Pr`��KଳcՓ�R�s�!��fU&�5�3q�dF�    IDAT=˩�A�=cE�V
��`��#p�9gᔓOP�l�����_���>��]�p�LV&a�F����ބcߴ���]�}��e���$�-�E��c�w�d�v�ڮ36@�˙3g�1�7&H��>@�!���v�?�l!��,�������̙ö��$��>87��ح�����CS��Th�'%ɶ)�򈛢�u{Ed��g�̺Kt 8�׈����J��uYϐ?r��g���5��S��F�'<r��(z`+Tŏ�yr}�>�Do3q{�N�H�K9�ZU�Ӧ���R<����s+�t�x��c�R��{DxfN"'�[%w"N\���8i�P��+��K�Oe��|e���`����n�_~m�"��y���x�gWa�e`�>�^�?޵5��)C�"�i5��]�v���d>�`�.\/�c��Z53?�T��umX�ͷ݂�z�?�,�'a��w�~�*,;
���l��P��p:�N��N��#>�1����?���*:�
UC1������xFL�ɗ� m������?�6u
f~��@C����7n�1��� c�#UQ��WQ�n-R���X&�l&�_���-ظq3B��c0r�4x^;�b�ϡVӑ�r5�"Y%�"�U׽�wPl��� ���}���r�jl '0����LJ<�E6m�x���a�R��������[n�۶�D��JeṾL��W����bڴ)x�{ލ9s����ǽ�>���Pd�����s��� ��8�kt���ʇ6zv�e�);�w95��,X���o|��hZdu�7�>����>8Kny�_^���muC�b�}�H��l�b�����^�I�à}�/�v�v34fl<�M#8rA�W�(�Ir�f�� }��m${���8��`B�U��ӧN���?S&O�R��k���~(��.�y�	R���gx����k4&�+��YOMV�b�+��C1f��mn@]K�Y������_�Fk+�s60~�gWb��Ϣ~��H;M��=䘉�}t̴��堵XBkjƾ�$��ȧ�y��jt���޻���0�b�[��oƮ��F�+�йaF�v��H -͒o�i�1��O� �o�	޶-(�*'O�����5����Cň�������;���;0c�$h�۲��-G�։io^m���a�[:|��_�s�/����!���	0:���5s����O&OVE��W���[ѹq=r2��� ���N��F$n�3��w�6��.N\���K!�]�8�2�<E�7��Z,b�#p�7���Oq_N����c���[�v�fx.��B8a7MC.C0W��0q�x�7�6m����BC�5����E:nl`�v	s�Lù�7�@c>k֬ݲn10�$�!�y���s���߿��.�SD_l�/���C_�`�V�M7-������a9e�Iم@t1�kQI,�R"�J{Ke�^�X��}��5�m�̦�-��]�c�Yvg� +kߣԨR���8�#.���*�J9�|tK�+Rc*@ʨ%L�:߻�2L�8Z��܋���/_ �%q7'e7�����(�2�� �T��3ʔa�%�ʔ�=�f���HWE[����Uo9���4�^����Ὰ3߼���������o|Z[=Қ��i!����S&�ɳp�G?�5�|
�cG�6��e�]X��3��=�O9X0�,��/�a��C��UTi%�~-z�f
�i31��W=�m�{3
���	�6w�|�?��<}���:����,uہL�kBÓObóOb�̹�����_B���^�@��E���A~�2��翠ZҔ�0�Z-S?��N:ظm6��+�տ����Ȱ[�t��l����D_Z����ǐ�}�A3qwG��đ� �X��pQ-ě��_~*Yv�m�N���~�G�;4�Bg��Iq�Д� vH��AxK�2A�reqD��ԑPx�d :n�K�(RE9��;sz���x���a��8���ӧ�Ɖ�c�׺�u�u��x������E]ty��o�8�{n��cv����ml���pt�K��r1}Cu����b��:����`�e2(͝�3��ŊJ�|(R�!�á��N]*┭�R;cp�Ծ@�	u�2�=j8~���a҄��d�+W�s_T N
̢��$7�}��$	h�Ɔ ��aN���^uM(�����R`�f��[p`��Jc�����Ӂ�G��λ����9����~ӱ�rҩ������z�hݼ�C�`����T�D1߁-+_@1���3?��	'��?=��W��E����Y��w�ܰM�5a<Ɵv
�G/�Z�� 6?t;2��67���:��{&�[����Pܸ����2���@S���+PY;�~�c�#���=�tS=�7nEK��
9��g o{/��r+ڟ�3���_��g�	��c�-�"�n=�T���36*�};Ƽ����E�3Ϣ��'ѱ~*�vT�L����<Sي�b����i�N\�؝�G�*�lE�b^i�e�8�ķ�o}Mʨԁ��S��w7܌/��@�k`���X��D�u�i�N1#����"�#�N�u���<�;�u��YCw&.q����)S���5�b>܁d�����_㵀b4�<���/����& n���kt�p�1;v��#v�WK�?��M�wS�C��GI-(ų�=c�^}�n����8/\���2����̫�B˩����2/�DJ	���sՀU����jǇl��p��#�M�'�Lg�"�:���ċ�Ǆ����_����K�z�y|�+&��D,�J��ɧR�;aZ�Nd6��;�"T ��U8%K�8��R>`QBb�/5�2KYK?N�4b-�@�;��(7���S1�=���ɧ����`46 c�(L��1l�\�y���ܙ~O��!̝w*����[���Pʤ0�[��
4?�N1���Y���?l���(���a)m�w�qv�I�Ӂ�߻u�aԂ3P����Yu�Y2i�I��ytۇ9a,�~�B��O\�#�kjp�נ}�:���Pٺ��C�ѡk8��L=���T�|�|+ZkG�/|	p�ش�V`�XN� ��:sc0���~����<�'~#��܅jǅE��83(�-�A�T"�o\g��S�AIC2V
锅��<���wJ�2G�%w.�o��-�y��& N&��F|��ě�"��rb&Uʇ�LDZ����|��K�։�ĝ���k�.ZZZp�%�`ӦM�g��~쵀�� Icƌ�R8��|��q2�R&ҏ�1ŀ/�"Q� ~� p u�.�,X���|�;I9u�?�z{|q�~v݃�;�[0Q�Qvڄ�{�#g����[qQwg�zޟ nE6�Ҽy���W�Ų��\zVvySR-?��ʩ��;RR�m���s�qtS�Ab�-��G�S�ͬ�_��M����u̘1EJ:+^Z�/}�"8^��[�m�Z�����s�t��0���P����QU8%sh�~�<�{� '%)�
А���j���5du�Rn��ܼY�����&b�3/c�c�@j�:��f)Sg�Bk���M��9�X�<�D`�+XqϽ�f�P;f3��|�����`��. ��8G�}���Ч��G��َ\u5Vnچ�l���ϫ������)㡧P��HM���}�Dl��v�o\�(!;i&}����]x�W�"[=3.�ŵ���?��b+���z'�|6���<X�������̟a��Ԅ�8����B'���JT��c�h���D
-v-�#&"�6o>孰��B��;��PSp�&�`�N���#�$+vQ8g����L���왉�S���uE���P���?���~�ۤ�����]+��oo4[و��vaX��2����Q@�:좦e���O��$�#��bǹ+7@@9�\(��x�bq�n�Ծ�ڡA�oUU�4����`.�N˸H`V~l18�w�q�4�xs���l�^�U���/c��S'��}�{�jD�lI8q}pBZnYr�Ϋ~���5���m��|��K#��Q��Q9R�U6�u��^?/�ƴ�Y��9���W�ɲ�@\`�Y��i�C�M�N���k�,�q%v�R2�K���ʠ�h�p�oG��L;eh��Hc���R��ljck���
Ю,u�]����Ϗ=
�bG��',q���� Nq�<�tZ��$����E��,zp�A�Q�p�;�!�4�����7�Y�	G���?0�MsQy����V<��c={�{���桇�R�
i�@��	U�Cљ� 5d��v�?�~h�ð��{�u�c,�F���~�A����.�;�������KX�:�̙31���6�;��'��:tlތ��S?�y�����+~�aUC1���6�³W.ƈ�dR9�N����V�>t`�x����i%�>�dkj�?=���܍L��aH6v�r!=cV5�b�����5�K�`�_�" nH����J��ǮI!Z�^��>p�Ń9�]��w����:B/D�K�$%P
!���?��U������7�.�8+U�3߆%�c�@��76���$�Q\Y9�0��C�l�A�H+Q��52�)�/%f�a��Ɔ�Ŧ�8q����E_�K.��i���� *dTG�<oh8�7-Q�q�����rׇ��A㚚���b���V^g�d2�.0���FUgv\�,ts��1P<ꨣ����+' �`#8H�o��ێ���_>0bgCm*T]tZʐRj�04���R$��O2q��Q\N}1g7w� ��K���h�R1=2F��A/�}h>�;G�����H���aC�w�g��QT�� ��R)�mqT(�B���E���mM���%���[ae���������"E�<�7I����͐&�vF$F&�~
p�;�tp�Q��3�Mw݂��n�	�}�0E���U+Q��}h{�%d���؍i��DHs��&����1�0G���3�TWb�e���vy껑��j����h^�����|ׅ���YC��9��8�=(��f��=��k�c§>Է�����5�P{���g��u7�
UmͰ�3�B)DKE%ƾ�}ȝ�U�l%�x����fT�� �;0���}xj)����;�r@�v<�˫��ף���!`S?�$�HM|M֍x��w��3qq/�B��rl  #0���`U��9�9�����$��:o���7��{�hR�ѮKY��q�U���W.��X���L#��
K�	ur�ʉ���˻S��Yl*��ىo�ۏ�_�~ckk�[YY����i����}��C@G�-z�A�_t�h�S"�,����\r����u���04���۱�n*���`aUU�(��S����]�3'�<�r��p�%��(Ϛ��h����1�<�c~t�UWQb$���>(Vo����v���8bg�Hją$qZq��8�Wi}��� k���7��ِ��"�Fi�l|��kМ�ӂ�rj��F5a� ����s���F�n{�d��QR�3�\Eg��A��T87i)�8o�}�cG�D� �ж7��S�����B�~�[Nef��B��@i��[��)��N	�,W=���[b9��)��c����B	Nb�[ނ��#Ѵ��۷C۹hkCβ�c���Y}��Cs���::�����UC��j�+30vlGk}���Sg 3b�!C���й�U�������O�:]�l��#`T��;P�IL{:��5Eڄ��U���G�ֶt�]��"��fP1�B�Ð��0~�L�Ln_��p_��z����m��;�#��C��I(���a�4mـ����8n��Op�[3I��x��xOy����S���x��m�҉K)[��<�5�n띧��K.��L�����V��/��o�zeBN�ث�س+����ҩi `cL}ߓ�_''� �~���a�V8�B@��2��@9qS��;5���[�n������|�����NH���G�w���ڵ�T�0F麞�,+4MSokk�躞�u=W2$mX�q�'[<W�x�? v _�@�Aлp��+��3�H�H`�:ͷ�r䶟����v�米��*�������j�2�J����/2�>��^+�ĭȦ$����AKJ�\f�4UN����	���φŉS��^D�~�7 ��X ��)�R��ʪ,���w���RTm7X4+w�����0%7D�Q� ���A����X�����e(�%X)}��������bN$'n76((���������I���� ;�%ׅ[tQid�>��YZGG�#��@k+@�Rh�@I�|	��Э���tC���	��Pe�������p��DGe�WB�Ӂ
�Dѳ��BK�[*�RtTT��в�M�;�9Ch)v ���������.l�BMjN���dE�,�;��itC�4���6��D�6tM�S9����BUCm�f��S�3(��AApÒ	BFQ�w�4�fΒ��aX4�������#��k�8��8���`�-��H[�hx8f�\���!C,����u��[�@-�X:��6�׊Fi���x-̅�g���!�����<�P@�(н&�SՕ�*�ک�d�Z[ۼ;��s^x���j��<�0��\.g�J%;^6��|mss������---Sǡ7�pM�h�[�����{�x�m�_�hя���Zf�7�.��8��o����xpX]�(�r�3"��4�ȉ�f��ȱ�;c!��".�z>��w�@@\���L
��Uר�T��� ��8)GT	��ٻJ��~��t/?�;G�*F�ҥ��P�Q:���1#���6�ƌ�y�v[ԭߴ?��O$S'n��Ԕt�54`Gs�p☉���*!eq��� ��d�w���KC�[����h�(!��|�{0��� q�*��7�Ү���e
�˚,�����s%nCg�S����!mڢ�/�k���~�CFs�tZd�-�S@ֶ84�zkJA�mA��KC�}����4��*ǁ�%6��I��}|����x%�o��e;&���R��"����&aV�R)xZ;k���vh"c���Q�1 ]�C��sĐR �Xj��]�!ˆ�pϕ���A�*�Ĳ�8g��Y� 5m�b�vZķ�Q���KXt�<�,�����ƛ~��V�A�5V�c�.��+�g��S(��2U�4yF�����k�m��L5�M.��Y��dM��2��#׿ N��yhnn�.]��/���� Y�ٺ��zj�3�<�[�.jkk����0G�^Q*����@dI�k��4�����o~�fۇk������(����5�b�/8�8�)
XN��/��b�w�n)ǯ� .m��L
�����5�N�a���F3��3�k�uŉ��~~&NfnTo�,Yz�ܵ��mr�vNѶ���>,����RA�S%S��<i~�=����V��_� u��%�-z�# j�m8t�]�L AK:���U�:p2A\�݋Ĉ�h����M1�Q��<��H�%�g����	��zR
�{:\���ӛ�Q��ch%E�;���4E�5�2�;E&��T�S�
���ȣ���>��\A�5�����/��H��)�﫫�n��=��#�e5d�Jغ��@�/���������Д2\[GrU9ivQe4e��{�Rl���"�hpUa�x)�K��ld$�SNEϤ�^�@e.�!�/��"Al�|�4K���L��U�2C�*���u2P������k���zO�|	�6|�P�ʪBb�es��GE�¿��|��_P�@�ep�}��{���M�@Vɧ�VJ<i	�-%��o>f�8��6k2�._���{ ;w�R�I�' ,���]ޝ�ƆQ9u����3'�4M��ԥK�.��o�p���9������Ν;G����aÆ#����������>��4�t��IE*d�Rm��Y����2�q�w�A�0���?��{�����@���^g���;T��_ӭ���~�u��e�5�b��-���E^܂�WcyD=��˕�qO�L�T�6A���NG�  TIDATY�����F*�萌g��,_Uٌ�X�5ֺ믳�z������ի���_q�,�K�Z�����Ȧ,y�s�a��w��ږ!�թ�&�;�^����J�tŪ��엿.�e�T��\���% ���d�LL6tQ]�㤑Cpz&Dm~O�8� ������8Gj��B|������~�2w*�jeI��ko���n���i�yWǣ�:`
����G*��"����Nu�7�j������غ���N���&ڶjR @e�v������N���v;��:��Cy�oN�o:Php�]��x���af�S����m9���E����������ē����fܞzf�	�X�Z�����	u&�È��`��x��ކ9�'�Ԡ���ҥ�q�w���U&�
E��9�j�̆>�̞����4�̜&�,�����zr�X���o�Ž=P��|���+V[�n]���&K��B�W�a۶4f��/��!��,��5oD�Wwx�-��T+'��x=�51u]o��o�&��(��:����)!����_=4��n$�S>�ozF��uu��lA��b6�78k������a���{�����}�?F�e#� � DY��x� T%i@��5� k�A����qF���	�b��n��I�x|���fN��K/Y�i�GK�ŗ����|M�B����g�ʶv=�#�r����j�����d-Yh��*�a����@��]��Q$���-�OD\���s����j�x:�i���<��]��$L��~���6X~��`�<�s�9�={��Czi���7`��5���1b&L���c�"�6ŝ�?��x�!�y�x����\/T|Y��ɢ�;=�1o�t��g��/܁�^���o��6����@���87�:�5�z���n��J�=�V��fKJ9����J�2�]�a�}=���{��bª%m�T�#gK&�.��Q .��I�@�m��̔~��	�zfA��-�L�hE1�R��F}K[��d������l���C̝9_t!fN+eӕ�7�/~˲2[�5��q,�z(��J�v
��P[h����|��Ai�r���@�<Xz��|N]�I�-qf��l61�vM���bEQG����Wh(>��]�pH�	�ٰ�w������QG͑�&ŶI�P�f��
��Qpݢ�/����<y�1���j�+3,>E�Iu�N�1�I� �ƜY�$�;�2q?]�����GZ��A�����"�{��_=<|W�f�\���8�څ��Ҋ��Fe� ��6�r]�M�Aq�q�)2�M)�7͗r�Z�D$$"'cdW!�v߇+���QN�Q܀��#��)��oR������|k�G�Ũ�x�{��F���z���vܼ�Q�'��OG%9�YU��ҡL�RXB6,��DW��3�>˩{͞a;��k;�T�>��*ǳ�ńk�鸧�ËN���C@ �֡#)ޫ�ADWL����Q��Ì����O������FK6Χ/mʘ6'�b�4Z��Іu�6�/�?����OlڰQ4��vy�6�k���ָ�:��ԳϖI�4��o�F>رDF��56?��rj�G��>�'Ĺ��y�~��YN�4����-h�����(N\���c8�M(N��U�7X0�ُ�`��.-�GJzq�-j�oA�������ٷ1����dn=�8�9�V �666�t(��2'��ǎ��v�|��W�q1�t8n	ͭ�q]ܫ "��0X.�@�R�/!���e�F�'���9����`��d�${F@5i��q,�|`Y���!�l��-���,6A�(�+$��8y��Nyͥ3���ٳgb޼��8a��Mkj�!�� ::<i ؼy3^^�2^Z�k6lDs{,�+���I'�Ai�]�j�.q���i̞E��.�Kʩ���Y��ष�p�Wq�õ��F�4���d�BI���&���)�J_� N:���\z#1һ�Vŉ��rچ# �h�د���ZZ)�|��I�[��'+�Ą�>c�6q` N�3f�,�G̲�ѫ��o��g��}c�!:T4�V������n\�⸕�( nX��G)N\�>�S�x'�(�(�*tɇ��kxms�C^m!E�T�8ϗ�����sai&tdT5 �����;x��ՇVV"e���r;v�d�≐��c@KcꛚaR�%�fCk��LF�2�aZv�#�d�t ���,^|�7���&;?�H��>y㒛go��G�l[A-+�J�����"�	JZXbS�E ��rz��Q�y���6V�m��ƙ�\�&��i��`9�ٶngJAA�!Uj��d�A{���p����9C&�E��-1q�$'�8ո��٦%$ӈ�$eA�i��	�(e�hN�@����qzh� �;("�����J'nx�Y=(�����@���$�K"0�#@jI�c׸��e�@e��
���@�j.�%+F�(�UUC��א�m�wq])�0��9)��wJ��� ޻�cei��3Mա.K���E}AZ?D�Ը�Jw�9��z���_4�Ozrp}���AHn�i�����#��V1�\�L�8ih(.��)M�@��
��%�B��@6$F6V�Z~�e�������>����u��O^��9e!0S� Bg3�h�'��:�[.��I��R"q5*� ��%��ム�8�&��B�� `ĥ�fCV����X�3uVDE�b���I���9Ê{J�Ш�@������9�\�&MI����H�0�E�-]�S� #-����#����&M9j���py_����x��Om����.���?�=ޯ�?�d��@�$����yR��(�����H̉h�K�,��%�|��7�u�8H@\���7LYs���^�m�Q���<hVŒ�0�@�-���%J	ď��q ҁ:X��C�$(P!*�
4����euZo]����/��b[p*-v��SD3HR2T�R
�2qĩN�����Q`�TbV�^��sn_z7��j���q�� o{v����ĺ��c{��	�,ݖ�86Cp�)������0�6q���nȽ�W����.9i��b"�d�o���<V::�B�9��)�R%ה�J�� ������73�~�H2)����Ш�hp�ќ̦L̜1�~�S"1b�;����Ɔ���Y�����Z���{o���7��}˶��P3u/�,;�:�g���k�����# "�47�>]4�cf�)¼�����?��kD��fK5��a�i�r��R��tfs���3q¶�x��]z\!\
p���G.��.��B���ʩ�E�*��qfP���%FK�\�%w-E}s��+�LZ��w�S�p,r�9�r#�Qş Γry@^����Jx Ʒ
zx[M%�I�8�U���&���)�.�]̾S'>z�%�����apā�������,V�&�7{x���CQ
�h�@+\��b�=�dRV"�]��]7���=��D:�F��Xr�k���ۑ��(z�����ł�����	�O�7�Q& ��k���Y46���r:
i]�����G�͡@��4�J/��\7Di�u��(���\*�>�h�y��~���� �&�����NRm�=�u��d�s�6|�=�=��Z��,�/!m�\�$�	�T��
�Q�I��s)W⏆�(ӨV�@���'���w-��K���� ���;�}��q��\��� �R��hY����F�]c)'��z�����*�f�0���� ����u���}����Z�^�{��r=e9����"1rw��%�Q�2q�$H<Ib>]x�2Y"����}�@�����we�<�h��I�Y,B~s�Kc��Y���s���Yӡ�V]��������_�ڵ��w�������K�!<��Q���u��L��#W�_)�ٯ��~��sCd�"g��~�ݴA @N�,�y�ݒ�k���)�⛺����{[ʭ���_AG��O���
'N2B>�uq$R���؉�pBmޕ0�ж𢡄�(����l~�/~���}�_u2�tFZ@���V�4ͬd��g,�W�R�-���PU\61���X�͛h:vw�Q�eF8��@0�[,CÜ�3p�Y�����Q]``��7��ֿ�Mr x��l=Ye�G`�/��������/|�K$��K�~)t�6-�C	����6{��r�������%�V�T�e��k!���߅?�y'��:���L݁-��8v�!s;&�?,��q�Mթ7eG޳>L7����c�38�BCmq� ���WPy`���D`�E����S���ڢ�?vxXYpQ�S�,]2�i>'A�E���!7�8%��cٗ�p�uU���Fl�W��i�x��VM�N�͙���:G9O<�_K�P�'\�Ňz���V7���a?��7N\�|�՟>��3�\��J�!,O54K8q:g���)c5��g&N�]��(s��ˬ4��L��Cx��G}���I���E�3HL>����VQ�"�;Ԑ��U���[J���M�l%-���}5a�i�TZ�t���Mvd/�q�| �.Yg F� �D�(�TC`�<�h��pI�5)T���a�v3ӭ��U(2���$�g���	�ys)���?�cb�05x��t�Ĥ�cq�'a���;b�C� ���\�Kվ���$π�y^�Q��z����x��S�-eXH���+��Ŏ���W0U&���1���S��	?/q�:o]\��S����L��*x:�@���ELtoK<C��۞	><Ԅ��`
��,�;�t_g��d�g_�a���bYz8:Ÿ"{p�<��|pqK�8`e��8�1l4Z��,)S�zS+
P��)�d���!���gO�A� vO���o/M0QWyWFN���U׻l��f�x�E�mK��h��Z�aq�%K~����sy�#I�+�t?/�];�����O|j�I�F;)��L�VD^�-˩�U��JR�Hڣ9q=A\7g-jl�E���'y����LE::20S?*.��y����5u�����a��3
|��`�<�j�6\w�S��0B����e�]���uc׆����ｷ7�K?ƅ��߼2��S(������4�bt?��!�HQ{��2�����C*�^B�n�%i�/+Ê�cď#?/m�~v�' m?c�aq��%K�H@� }���J@�!�`��+6̿��{����>~4�j�|�V#W��(��줨��w�|S��owjy�c��׊{y����O��o����6.���uO�t?0�(c�=�����{��N�띨v�C7^՜Dɘ�pul*`v���u�.+�vwk��;G�k��߻�����/?�� ��m�V���ۯ��˾ݗ�O�5�#�������]�v�}�?��s�9g��X�f�?����r*Y�$H"�D`�E� ������;���o~���L�F q�4��6n�x�]˯9������UUUR~�g��Rh�9�Ùa�$I[�iJصkW3%F.��ҟ��';H@܀8�w�6m}�K�������a5��y4p4�ff.Y�$H"�D`�E�-e�]__������ŋ7��29�C�����m?����n�����N[�j��*u]7,��� tC]s�0dg@��k��{���$���������n��Eav{aR�Dd3$�o;����:l��`����tI�����|Uۥ_<�~=�{�����A�S��z)�F�g�>?�sѶ%F
�����>�=P[z�����ǯ���ԇ�?ߵ�8>��g_Z��.��g����6�9�_syo��X��$�)?�����6{�~���������9���kŽ�o=�K���\�/?���Z���'~������7���,���ޮ����������b���ӑ�x�$�Ƃ����}���s��/����{�y���j<�_���cǥh�
�1*~-��m�5������gj�P����%�������k��Ѻ���u��"��,�ð�T*mhjj�z����7�E�����sקG�!��w����}z�ƒ$H"�/�pg�����Z_�n�>u�T�`���_,t��݇�O�$I�$H"�D �@��$7�OPrxI�$H"�D �@��E q�u�D �@�$I�$�H@� <i�!'H"�D �@�$I�\I�$H"�D �@�A���r�$I�$H"�D q�5�D �@�$I�$�H@� <i�!'H"�D �@�$I�\I�$H"�D �@�A���r�$I�$H"�D q�5�D �@�$I�$���웙�����    IEND�B`�PK
     ��/Zִ$�� � /   images/4fd5fc97-bc4f-4740-9bc3-7af0136a9299.png�PNG

   IHDR  q   �   ���d   	pHYs  �  ��+  ��IDATx��W�\Wz&��kӕC��aOO6]��%�LkF+M�hWڈ�]�"vc6�i^���;��X�c4R�gZ�ک�d7m�M� H��!|��Ks����Ͻ�Y�* $ �
u>2q�2o^���o�߃��������Œ�%qK��YXXXXXXX,AXgaaaaaaa�aI����������%qK��YXXXXXXX,AXgaaaaaaa�aI����������%qK��YXXXXXXX,AXgaaaaaaa�aI����������%qK��YXXXXXXX,AXgaaaaaaa�aI����������%qK��YXXXXXXX,AXgaaaaaaa�aI����������%qK��YXXXXXXX,AXgaaaaaaa�aI����������%qK��Y�o��o�A��$��QJU���y�C �ϴF��N黜�-��车��B�G�l�?S����YO���\@�y�e)���0xf]���v�Uqr\�q�.yI��y��r�t��:��o�����������F���r��;EG�%BF������Wyn�5��׹���=�������W탮�B�g\}-�^_>���i0��e��1��h���ޛ��>���O���0�!�������u�ǢHK�k����&|����}��'z������s�s���/4���˜�7�U��ՠ��"j״����t^�o^t��{�,���_�ӣ�O_�0���:��8�9��[��ַ�a��`I�2�;�������������Al�}��$�K�wVԡ��ZI�jβ���&cR8�o�&,�a����@_��ݧ�o��,H?�5�u���g�1���|����d��\��ᶐ�}�پ3��#�s�knS�w�Zg�s���Z�(�g�7�ws�� ��7��XG�mG�g�k�l��Vk�������=}��bY���e�j5��X�r��_���,˺�:P�@��<"����&n[�0߀`aaa��p]�D	Gi��푋/�=~��
X,;X�̑�����-��F��O/&p��Keaaaaq�Ȳar?]����eK�9�<�Q4Ҏ#��KB�8��3u�|���v]�����s�,�,�[���O3������H,q���D���wx}�������3�PA]��������12�����98M�ásX�l�<�Ͽ�D�ܼO����v��U��������k3�U��n���o��k��\�� ����|a�: �n&sE�2�%qȒ�Q��K݂C/&ti�Ηd����U�D�*���\�r>��rъba�~��9��Ƨ?{�\$�v
3���ICN�@FC��g�KRI4uFD�[$��N�υ}]"�-�X��6�:4��3�i���4�$���9|�P�̤-i���]y�{�#�v�	��zw?J������'��t��o�gtpiD.���IDKϑv�S3�U&�����c,݋X�|�}��gc_�!,�[�\�a�-o�I�%�H�����W򟅺L���Ӎ�j�x���)u̎+�FF���ٸ��s�Ş�"��Yx�!΅�L��'�!�Jiف']�jf~=�ZX,&q�l<f"Y.3�Bt{�ͰUN��=u�FP�1�^$�)>���&UR6���N���sk.~W4A?�#ɨ_�J�t�i� �	X1	�;����S����-n,�[���$g��I�$p��ߥ{u���C��Ӎ�3>x�|S�m�a:Ϯ��k#/\��;w�.>3n ?'���%�"���#ҘE�l���I-p Ifm����An^ʒ>��C��}9���~�8E�3�X��Z9q�f�vT/��O�.[�5y��<8F�~�K��@
C݌E>��~Lm�I [�%ً��jl�<� ֮���m�N��(e;��K�9�0l��K���r�C���	$��Q�N�'���G������P	k�s�Y���q���!��
���^�,��̧� kc�Uxd���P�Q���O�{���R�2v[�~�|i�0��P;C��K�n�ı�LbI�~V�R���jnT)��|��Y��g���W��#-qy�ߪ��R�ұ�)��ލM�6aӆ��h�X�����%q�o��F�^�W=�U�(��Z�v����U�/���}�¼"^,��'��w:��:�tff&�.]��MOO�g�yFz��������#f$v��7]Z�:��1�,���\ܛJ,s}���=�Awcp�Y��f�[�xBɭ�LK��)��iT�����5k������!,,�&r���:wԘ��)��-�>}��1:�p���c֘p���2�e�4tS�L���cP���V#_�/)4ӟ��ȶ8;_�Ln�Zܮlu�8�L[�dq�aI�-���㡿�����&&&���x��NK�s4��0U������{N���Ht�|���e\6��YD���ğ��6�}D$gh͚ջJ��č���[�g铄�;k����7�����o�g1yJ�I�gb]��Ф4�]b��wQMCPqPA6�0�[�ڜ��ma�Ԡx��S$ڐ��QR�@��>����b�8���gE웙*�
}.Ӓ�)�I�퐓�T��f���9S�\rc�0GWڤ��y�����)BOa�ؿ��Rk����LMM���599�xI�J��dN��獹YS�� ���$�[���k
�H��p,\��R�\ף�}�}	J�x��V9����kfx^�i��E�u�j�fW�#���Y���<d�\�����g��L��.���N��A,,>5���"�>'�F�P;hQ�iS#�~	q#t�n�!�B�a*${�6R��t3ů�a�1�ʌTHD[�p��r� �Y�#���r�XJ1��1���p���MlX��$��mH�g�R�H#���_�%�2�����k]�͉�9�1���;(&sL���[����ZΉ�Q��Sip�v>_v����)i���|���������{ڏNh�b9�ܡ%��]ޟ^rE�  a9�FK��=�X�p�Sې	O ��9D���HuUy��i������)K9;B��r]X�sU�*m27zr���u��b�fȠ�E�uK7�6@�3�;��2���%���&r�nb��԰$����ñp�v{aZ����ۺr��C�Q��T�O}�����b����H�$7����Kwi�^�����P����N1HOeEPuq}��aɛ�G��(4����Nsq��$�ݧb��8S��"�'�XД�ɩ���4�4$�7�"�x"jb|�4��t��6�m���ź(ڱ��w]�;���<�5ֿ��봡y�}���%m�g�ٿo�m��r�%q� �D �%�[��������d�}<���@��T.���q-�6���lكO�2>�.�r�,I p�6�겒�D�v����P�ɪa*(���Q�r�"+�ڨV������H'1�򨛞��$"W�u��N�������[��p>V�֋*���f���K�n��0bGws+5,�V�ܷ�}K�M�S�����o��~D���hǕ�$���&qE6����.��R���+3�"��1W����_��ل��?^VZ�4$\�>M�h�q�*�b�;�4��$h�Ho��[88��3Mu�,�PE��?�*#�f9n����ҝ�x,�&���-GXw��T �-R0��ԭ���г�m��UN,q(ñ{�^���x3��^�����xX�P��˥�H�LM���&m�H:0ϸi+ni8+bޒ$�[۸Vū`fjCuY/Oc��F�{���BX���X&}󉙗mK�eq�Z��-�,��(,q����do��fY��J��£�ܞ�j��]^&�ڑ�$9�.�c+����.�4�܋�9f�v�i��ocKt�P{��O��	�Y[K�[�1uf���נ��\<ԫ����}{�H\2Ǣv����o���l��`Y8�;��S�yn�z��qaq�k�[��$���;mz��Ģ����M��;7A����Ȅ��sH�c���#p�o��K����.��S�vi�Kd�`;X�a]�&��U�k箬'i��9�.���Xï�,VI�ª�aܷk��^Y�o��|�q|�o��T#�Ti��a%�
gN-�g���r{�6��b>	��o�����ÇkD�r��[�e+*���c�ِ�K��|Ͽ-߳�*/�ŉ��g�g���������B�����*S�|��ַ�uk���bXw��M�^��i?�`��q->+����:r�S�"Uo��[��}��A�s���Sඓ:��P��6��]���gZ�2�����80'=��-���D�b0���c�b�uҲ�%,L�b�Νx���Ɓw%�N�F�w���?0��X�M����E1��. ��|�;��߿���_����G��Lވ�y�ވd�L��XQaD)o��]��2W�[�z��3����_K֒n�*'�~���������Y,����&[Ue'n�_�:t���ۻv�	,�H�%pK�����U�*,`�Lv8��T�L�)Wba��<OQ�x\��<� �Hc����00Zt�j��߇����GυZ�f9�I6*f[�gO���Ȋ�W颴��9���矿祗^�*a��D�6:���^�c���$��X�o�6ew�|�.7jSYH������v{��E��G���,��XJF���xn������F�M��!��}j
՝��m3�,�*>��F �E>%������}�فz�u&ք�֍�OD��\ײ|w��Z����f��l���ߔ#qg���������q
U7U�=��C|���޻�6oD�3�S2/�n���=�j.���S����.]��TfgZ����JgM�TA���z/	M��sp��zD4B�`>]�B�|�������Ɗp��8������j�����T{�ȑC�:��?��?�B��:�kǨ�`��R*f!0��]��xkD�^x�~�R,2Xgq�Ô��lp=����)E3A���iZTmԾ�a�xiJ)_84k�R�ф�� �K�$�w�����3�?��V����WqfR���f�r��U")��=�qO<�V�Z	n��T�@����i������^F%�\��{���(���?��L��l+f�P��Pq�J��B;VQ[�t��n�7�t0:j�uj���S��8}�^��E��%����B�|VU�W���?��[��������ĕ�z�ZG��eA�^�V�$���y�\
�����o�g�(+�zw�� ,��X֐ؖ�RW}�j<��+_~{w��=wm<K̹t�of���6���+|r�Tf�E}����j�\�ՙF�O1�zv�ہ�P��y��x[wn���Q0)]9����^z�U$�)5�E��*qcX��(�U)�u���'�g��Ŀ���5��Tu�_��R;Ȝ
P/�4'w��x�v� |�����/�\��QᲐu�z}�����*��-�g^*��mƫ�>w:޹�O�<��/�wb=�I.4{�?���Ѳ��4�7>o�ﳏXZw7�ȄY:>TA�]V:V�ab�4����ޏ_���&&F���'���hyi���������)%H���p�����86��FK��Uy.�o�>�Z�����R#���{N��?��&=�<�ܵ�lZ��|,�Q�l{T�<Y�������?���Qu�R{6U�L<��p����w1[73"P��� �Sg����)W�\���0@�����â̱X��'�"|"tY,�eI�L�C�mI&9���g�Y�1.��Y,s82��uI�z3l!m�I:E�5�,��W\4���2�5�8KMc�9N��h��YԾ'Z��7�S���3��86��S�ؽk֭����p��q��y���;DvB"vV�X��~t�K�J��j\�Z���w
��C�I..��n3ưvP��8^,q�>�5Cڈ�*���%�3���լL�VFT"�Kd��r�rQ���ިcRe`�}G����>���z��R�T�|��!��w86X�SH\��/,JC�%q���[� �\2UJ
���҈���r����p�Me�Q����K �ޑ]���uݩ�ᰰ�Šv��ݞ����s�n4*�n[{��W03����8��1�ۻ�z���?��?�J�i��BN⟮�k�Hl2� #ғ钂j��E�e�yb),.׎�o}bZ�?��2�/1��:)i&!$7���i�F������w�y��ߨ?�Ui��	j&f��JG&�ܿ����M�D���|'H�\�_A�k����s0�Œ�)J?�w/_�k�x��u���/4u�y��B�_��tSS�f&����d�"�)%a�k@r͕'!��܇�vH�GM����ً�!�4�D��?z{����B��m��b罻���onٞ�M�W�_N��~�X�e��t��$`i�}R�8��Ɉ�9�k3�g.17/��:N*�\?�T�х5�Ɨl�c˞ID�^�1��.̀�s7U���zu����OX�<N%�!�#x�q��䍉9�WyB�.�ۉ��W]��G�Ud�->Xw�`+6,=t3�ʨ��d@!�I�V'�K������I�gf����s�3���s�t���Η�t'ܡj)���C]��7�i���5k��݋�+�	5O8}�,N�>������^z�����Ѩ�$ku��1<��}�O$N���Ļ�j�J"����Fy\��H�3YrX�%-�����s2G��5%"y.�ey�
����~MK�4�.咊gwf�?�y�IB4����2K��ρ�g�TzA��I]A0���\Xw�@�����7����ӿ���h"{�5x����J�
~�>/��2��'f8n���D��\ex�)��I�/jKV�<"R�^<�������o{Ej?,�/�O�đĽEI����f5�F%����u�6p�>Ǳ�?�<&&&��Wtx����+_�������;wbӆ����)���#O�X@Xy��,�'��(t�8���Gdʍ�A@�á���<�|�c&��%�t�&�R��J�O�d�rS�z:G!&&�HJ�Q�h��:���$1��L�,b�����/-��ۅ���|�T^�+E`��[ �N�2����*D~���z��L���l��t:]"��w���~����E����Ґw	��R�=�,S�G�k�Ü����^i�V,K�,�Ci�ap�T���<��jNaϞ�ر}�41n�U���}X�v-Zԯ��5t�)lٺ	"��+o���غm�$>t��HEE�\���~�E,&]NLd�IǨ�t7���&���r���%+K�XɬUIF/����W���e.�l3�X�yY�,7�
v��	�v�(1�<�q\WC!D��u��X:��y����#\���r-Xw��ג$qK��9H���w�خ��������Aevc9�������P�˗�Y��N]d8I�{��y��dpiխ�(�*>#nw�,���)}T�������$�=��ƽ�6�Q��0t�;C�`���Pڱ�+DI���H�6-������k��ޭ����h����'m!�k?����=:��e����
�3�D)p���85VH�eRJ���$�����S����7�T)]�D,�>
m�e�EKӥ=q���0�:^[�h|�!2"�\٦$qs���4��ĉ�!,��5Ȉ5���`�d�-r"��ٙ��,��Z��a��$����F��W!�kJ�tk-ZU��)w��-;�����Z|Z���-*���g�Xn56m\�;�ʄJ9��IĂ�������k3Eh�uq�eD��\D.�UWw�؁��Vaj�%~Xv�>��(v���k1�Dp\7���Sq��<�QK2ٞ��*��N.��\L�Y,q����|���A��Aˈc�}_j����%��ƙv
7m	f������v���SK�;u1�MeXw@�$u2�qc�5�YSRO��5}��9�A�n�>������O�|�������!+�����UiR��H2��X�i��V�����$n�����0�\���&�M:t�aj�-�ӻ�}���{#O��������hK�,�3�4�WAq=O,7�7�oڴ	�v�(�9�2�I.D���B�p�$�Q�*E�k�;wb۶m8~�,�7i�~��񰘑�D\�Q���&��''8h���J�83Ո��:�t�����§\��Y΄k��H/˅�>��)g�ґ�T�N+�C��k�歈ȹ����4i�7��>�F�SKܝ7. K�n�o�~�g��߈5ح��)MMZ9^�:Ūϼ��rY|���%-~ϟ��~�+�9��r�����q8���*H��e�>����5������tlL�f�.�Avn���<6�K���j~[����j9L,n���~�|�+�r�]���{ <e��*�Sx�7��{G�l�򉸸� ��V��C�x��}xp�>!4+F���{��ko�Rld��b����r˸]��o���~[;�J�P����hBNPe����If����Y�9wO]?�8��F����h��'�pxJ!��n�i#DK��b���v�%ψ���Z������ǐ�N�"�%q� �>�([�^�ġC���?A�s���ժ2���.�G��1�v*�R��L8�tMk�k���,���t�]�?n�T�	sS�������|VL�?�T]��Oe�֭x�'��U�:&��������_$B7@�V�}*�	׃�Po�b���_�vn��aW�}�݇^ƕ���gw�X�`;!'�wR��0�90��=�&L��ja�q�1y�O��6����u��U�b�L�bn�+���נ�*z�N5q[ڀ�D�t���i�y%��y���6��.1E7��馺����q'I�r�s6�\����`�BiY�/&��r�^Í*�%\�u����-�"m��lU�=�7��rJ>�7&t�p����K}�FA�x�"�T���~b���J�g������+\1��L-�|���~�l�m{��U��67]	N���U�Z������wIݘ���w)e	ho�*�ou��A��Q檤������ő�$����H���(�{,oPhs���2pV��NB�=ݮ9�4�p���Jhq���~]*s}��[��t��͢{�;��5ty1i\�(��8��9���61�&e}U|�ϻ9�Y�r5��c��.�Y>g\2��U�u�]w[yq~}�Py��ޮrq�$IE�A�k�)�P,h�.y'��x��p��8����zە� :�Ɉ�iN���Op~|���c�k�=ز}�?r�NG�:�m+}_�`ڕ[�Oi�;,q����e3#�_���垉G������eQ������Qj������zzk�T�X��ȉ+�i��W���}��|�ݩ��i�.�4eK�9�!]׭��-�$7�R.e9��q�;�*���$՗ֻ�@'�"��LE�L�}�zG��{%��Ոg�5�͋c���3U�c��i��"�BK��B���	��E��\If_1Ҍ�q�<hԫ���p&YJa��4�<F��@s��Z�`<�����\>6�ТM{4�瘖�S�h�!uq"JǑD)*y~r�\���Z����9&��P<�#�G�k��XA�هt⎇�������U,Z�I�_�����q�O���H��!]�ܐP)	D�W2G���,G�-<���-��ڳ��!ۉ���ʳD2�<���}�)��|AX�T�+5����Re��N#B@���u��Mڠ[	�D��Z'$�w�� �meQN��::p��g
�Z}ڗ��Mς����g�148"כ���|�D\��}���@v:L!ج�/O�c���Ni��w� M�QL��hw��@���o7g��X�˰��>ؖy��O:8�b�
����d�8�Cڲq�z�)pЊϙ��<���8s~��5D;�e���M�`�v�#�jgϞ�/��_���y&������/~��\G��45��k{��s�ɳTD2�N�?����9�	z��3��c�޽����_��_pp0��C|<z0[��������{�?���ٳ�ѽ�H�j��nג���g� ؟l�����A�w�y�ݎ�HaI�2M0�,�Y��D�i5����̲y̲Pt;�:s���=��rd4F�X2諭&b������^����6��6uସ��ƹ�q�檷-!/I*��pJ?����6�zz��z���Ff�-���:V��G"Qi`�u4�hp��r g&#4'��Wk���}��`�!�	�d2AtƐV&n����ye4�p'�i��oT�Dy��<y�1A���C���+��[M��J�6*l�c
��rϤ��E��.!�&�Q�%މ��$�I�+���-U��r�G��D�3��Ę"���j�vk�#�5�5OHe֎�Ķ��%tn	ݫ��Q!����������J|�yR�d!&�����&ߣ��jѵ��w�5�H�1�w>�D֜�[�AchM:�
7n�L�gffPmT����2l�A��v+(cY���G�0�3)�痎q���B�N�$2��� �`�ћA���J ��!�LΆ��er��ro.���?>��N$-G��!)�Ar�F��<H-㋗'@�o��G�#�09�k�_B��!�r�ܶt1+�}U9�rԇ�<����f<�Y��ַ�u�_���7�xc͡C�6}��'L�����E����!r:D�2(�u���7��/оc:��D.��"�%q��Kqǻ�;�y���������/���2�}����6Q�����f�TZ�	�̴R����ހ)��E�[zGHf��&.��)�i�O��D��h�k]�1��]�:u��)�؞56���[QY�
�k��V���D#�8���W0}��=�Щb��Vs\�D�"�Y�n!W9�
�f���r����BӠ�B����bh�fTW�B0<�£��׾Cvz�H��N�NG��YDg.b���B��q�o��#�~���XROKI���gLb�N�a��c��c-�'G����8��Md���3���[�`t�F`t5�U+�5��u�[D&fp��8fΜA��qD�/�'��'�] .J�1̺Df�T�>|��i"�3D�F�܃���ݵkP[5��+隚ڽ1��ԙh�=���Op��98�X�q5�X,�l�c��WhL�N��e��z�b�W̵<��_�=[�즬��-{y��\��C`|���6��b�m�]�n�t��q�����+p��$�0=�ı'�JW�6�^��-�b���5a2ء��[�A� ���d�';g�~�iҕ��}�ex,��מ�d�M
������w�����G��:}���K�.m��G�\}vm�5��r�_O�H��fk�D��
x^=U6��UDp��󃝰����3p����Z�e,RX����m��`q]�RYp%�Os�uN�����ge�U?[<\�seD�\��z�~�ѧ1Hoa~)�zƍ�-���y��?���}O�&��"ο|uv����<�[\cq�F�{�I�<�0�j04@$���L�[�X�V�<��o���ob��9�ֆQ��nN�	�ѧ�m瞱��OT��+q9��"bS%"�r�v�ؽ�F"Gck�A�g��c�L�����*�+Y[5~��eSo���ﾋ��E�}2���c�%�iJğE��A����5�&Ə�An��Jo�=:�~��8�j��i�޳kzر���5FÂ��h�H��(]�щ+H�z��ڏ��Ï*�
݂6r:q�k#����D�32��]��r�T�X���L�b˒��m\k�}��D��/q��_�:'19N�.�DZ��S..��۴�,�k���Y2�7	����k�X����;��ďK��PМ@0�*���s8�iS��e���u�-�;cY�A?��O ^kO��d_<sKJ痸��E�q9*��K����W_+&)*t�l���J+��ןu�5��Bϕ��~����&�%�u�^��Ye�O��OԞ={ԕ+W�����}s�ժj��N�*�"y��^J��j�f����~p�5�Kv�NNN�J%K�}�����^�b�%q��E�B�e��l{\��]m�ӳ��?�2����:*���P��qXN�Y\E��V4��z+F������o@�m���ĥwX���I&}�D�}�W%rŖ2O�,S'C[�b�+�"x�i"o#��J��(�� ��D�F�ذ[7n�����G�b4�$��a�k��c�\��M,"�Y��E�|�D6�v���ӏa�>"Ec8J���3���2�|�ux��2���ٸ����bh�\~� .:���"{�h��n.���b%.V&��8/n^mR/D�٤���m��~S�b����l��g����� ��D�����"/H4��r\�j ��kVa㆕8�B�K�|>�O.�͡K:�������������/�����p�icF�J��*�����[��wq�'?%�5�AZ/�LK���2i+�o�ZV��߄�,"/m:��hr��a3o�\ek�b��Ko���]Fז�|\���*,��#�2�.�
�'/v�w:�$!��j=�C��UO��1��y�q��%�l�D�<?(�pM#�JXB�0�]��8�#m�" r��թ�>,��>-��]CZo��-s��+��p��v�=;ޭ+\f�*c��Lj#�sȖV�L�g��b&��!"����h���-�XrUr9U�`��}_Z�faN$b	C�VM-J�Ċs����pC����)z�XM�]B�B�sa��!�Y���\��W��}�
>y�9\y� �V8�L����9i��	�g%�f�C7����}�A��]�΋���Y ��y|��W�u��5̋s�˭�ҹ��MPk�`��M�q��W0��GН&�l�c+�gn>f&��JcQ�#�{S�%�?gM+/�$����M4��20J����z.��n=ǒ)LٝI��o��]<��,@������>�:>�6ݜ	"��~�$b�=�|G�IQ�-SBȔ���|���!���������K�6���5�����eZf�J�&��#�49 �Dn|�q�w(�A�n�Wb٥sٲ+��3��d2!�,4q;�1�H:�"S�CM�<WUp�U� �3I`q���+�?�ox&rR��ח�L-Y���M�����e����F��l����zY��"�(�>�Y�nX��!��ĩ��Pg�r�^�L�v��!��G��D[)��ٚ\R�3P�̰�R�]�߹��Mr����*V�L�WL�R��I�|&�0�A.I�Ӏ�U̸{ x�"p�2��E����[�R }1BG�C$f��6�}��5��`�,&Ϝ���K��$M$��(���u+����� FV w��3GVW�l�tL�G�Ό������Di��9�X�d&Fc�Գ��u+V���O� hN�`#����l�r9�Sx�1$�1f|!Sm"��|�i4��*]��H�y[�Nֲ0�ԧ����̱E��+����jf]����p8a�YH��M�ux�6�����%�9c/�]�i���Մ����h�[Z{�z��ѯ?���'0s�}�
隴Z�ce�0��.�"c�����@�s��޶ΖMr�8�Qj;�ȹ]׫ݹ�G"��qk��B�&&V�?#U�φ;���lZ���b��9DHc�n�u�<S��M� ��'��B�L<��ɯm%\L(��d|�e�<�,sw�g�ʻzk���EG�77�;�Ɋ,�lz:c&~�]C>�0ED�-ܣ̥rm,Uf\�ت.�3�F��CW,�~��*�bL8����Ȣ0����i����uk��H"��\&��6y��P�
*#C�AE\�,eQak_�&�1jw�ҙ��zY���[<�6�X��a�{�a��oÈ�,��pb ����_YarkMK<�S�R���*��'O+c"R���1(F:/��v�����η������N#_KcwVb-�_���Y�����_&���%�X��_�u`p]Oz̀��c���E��i4[�Ae�fZw%|/ ��.����~�������FD�|q	f�6=��~�P����g��qv�.�s�,ړMV��n\g��\�-�Lf�T����ŧ��G�Q�@~"r	]os>jV6�2��D��Є`����}��u̷��t�X�gGgD��]�={�_y�5ũ{��(E`}�2VƊ��N\aq����3V9��ȕ2<��Jt/�waX%2o\�>[=���W��^�Z�b���#�mI�2�%q��%n�tI��a��)1'Q��L`����P-D+��P�Q4�D*^������[�����7y�.Y���]"E�02� �:BȣJ4���;��JYԡA�Z����11e�������|B;K��!f:*��6n����&�$�x�Σ����p�==Tîg���� ��"qb4��ѿ�+4�;�9�4����䩐���	,��3��%"p���
�{'?�6���G0��0y��	9���L[Z����]{�����;�V+�3��DFb���7V k��͛q��I"Ĵ�@�u��U��Y�ӂ�8�3.TSJM���t�ܬݹ[cb	�5)�ĤD���_���?D;�D�9��H�Ƚ�����m'&��X��eOۇC%"�&��Iף�q�;���E_�)q�	1�O����{م��t�<����[��kO x�A:�A����*��'����~���1�ݣ�����kb�8NN��Ƃu�����O=!��eK'�(CxY�/7i�������|��V�$ՠk	��Ǎ�����t[�/#R&��+���Yu
�(ۧ4��x���d_V���Uy���s�KN&��k$y���ř��:�Ų�%qEX��|�N��dɂ�"�J$�-A`2�-�D�bA�`u(9��lk��͹�&2�+I,V��OJV���7��9R�#rG�X,V�~��gp��Wq��w0@Ǔ�&��.��J֦d�����&�ԈDt�\��F֘LHq-:�deJ%���8����9����9~y�6��k��u8�6 �� G�l\:�1�8	���`��
L��9a�C����!|�Q`t����t�"�L�'�9��?�.���i1]������L8@�����p�א�?�}�{vÍ��53 ������8s� ��Kġ�$bN�ƕ��>[rX7�I�J���l�H���jظz-��:mץkZ�"c���}��� }�j�.ǈ]�qej���U���3�����A87��}Y.%!���U46oV�I�p&�L��L�Ξ�/��/�8?�j;������L�7�-�CP�#��nR����;<�5�>D|�cD��nF�Lu#����_���k��OJ"��4�%����L�{��o���`���믣�� q,�r�����d�֠M���<]�K�Yq�M����YX̃r0��v���AʵeY��ީ�)��XH�[��Y�+8��_~�����r�dוd�oL��\\��6¿NI�
���c��jB��f�t�:��������A�{c�	��N�٨�Ț�Xw8ɲɖ&��0�cόc��h��#��H�i�
�hOL!��k�����8�_~�����	�^�:�g/_&�X�"疆ã��(��[�DCZ�(�D�O��A���շ�9�ƈiU�\�uOH[���]��Uc�5��<�f��x�O�l���a�W���D^�������.�0o��JL�$�6A�#��2U4�w����%}73M��-��L�@d-�{�}�Z����h�Ȩ��c���?1�I.�T��>���Xs�]��<E�hl���x�z#��$�����tTb9��-�:��\����[G�t#��TP�G`��=�=)5U� ɶ-*yh�[��hƹ|����/I�'�t�,�]�ug�+�V�	�d��1�j-��Hb7%�w���:ͮ+�z���B���{�c�]��������2xs����eK�,,D^d�O?�$u���~\�p�o�@u�J6"[�؂��c�+Ԭ;U��oY[��^hv�ӑZ�ڸoz�#ya�ӽ����%�B��8�Ǖ8��7¥������U�#�*SR��]S^�q�� �����r|"�T�n��'�����6.�Aή�2�c��b"��v�� gZW�qq}�k�I�@H��ݶ��ݒ����+���� N���g�&���Z�i4�&�z(�rr=!C!�〯R�#��?��D���������c��]>�w�LJ"ؾ+��I�ט��\�0)��M�2W�K����1y�=8t/[鴔��W��]���,$�JG��mv���~�ڀ�
.X gS�;v�2|��\���b��!`�*z���3qE���>z�e���Uk�d����>�CGb�ο�.����։lU���X�FW­աi��Ӹ.�~���b�_ۭ`h�v`�zfkB�sv�sx�	LN71�e�)�,V�3����<����$B�$�v>�魯{9�^��-��9�]�����\@ng������Xv�$��b^�:���6n��~�B���/��E����ɓ��C�)g�T��<��F$�k��$�5�L� ����#�L��a���('C8��Ͻu�2�ڤ,��J�����M$�mq����˅؅ElˎH�_�c�I�ظ�6Kyek�����E�LOb��_b��9��g.g'�>�ku��:��T�T���K���0�q_��##��5�#f��N��������dD.+ZI[��(9�^EܙL�;t�E��1�.L:X����+8y��8�;9W��r��&f���I�u�ݩ��"fЬ�s���5������Ys��� �t$�հ��ul�$��D�3$a�{�akɉƞOį�P�1�<��u:������Hv.��ǣ9�L\Bvq��g��o�3t9_:�]���g�O��ټ�ȬU����$#�k��\����<�.R7
"��\\&��ȣ�q�x��������6��}�3'Ncl�+P��E�w%�w�#�!}�yt�t��$�~7�d�:���s6����x�:sȚ�녵�Y��j�X�-h.�l��`I�2�2ꉋp^�8���'&��ı�p���m������z�1�߿���?�ԙ�h6�����$�������Se�B�o&_Z�d!�p�������I�F�-/�Zs)$�#R!��	��h4h���qs�3g�L2
m	��0��D�4��shGa��ċ?����1�i3f̐�V�Dmӽ��w�).��8��~��y3MTS.v��OJ�N|̴�h�����㬅p��{6I�%��D3��[����7��1B�MD��fU�TUry�Q��H�L\�p\��B���ia��d3hM}(�_U�D� �8��<wi �ED8M��#u`�u-cUA�$��>�RS�l��U��|�tLm�Z!b���=�`�`��7b���c�\.-�1n��˄��1�;|nьE���8�z��7g�A	T;7�>r:�j�f
�7��+�"���d�����d�:t�Y������5?�!��g��N�T�ЅaD�LW��z�!#W%�Y+�`]8���oa��Y�׮D�ɧ��Wz�~���ދ����$��n���x�m�v�*�\e<]����e]�p�k,� bK�',�[�p���3�胸Dk5���x��w���W��
v���_�S_�
~����/����E{26�|x0�0�����R!��=���!cM9.q̒��C0�6مl�J]��8^�g����:�} #VI� ��#�$䊶�.ZY����&?8�ɣ�pv������<�.�� ����bIի�h#+6`��_G2X�"{L��4H_���ʊ��nD��m@GD�<O�ʝ�C}�:�WJ�-����'}�f���@�����׈��$��6��M�r�o�ft�Z��@�w���5N"o�֟�>'H�Y��q"��G�[��1�)
�'Llح�A����'�%�ȼry��_����6�?�l���܎`�(�k�!��5�$���Q������~L�>E:GH�oqV%gK1SERi�|̧/�Bפ�fF�Id��yH�"�k��b��ɋtZ�
�D�'�V14���Tb&RD+���������""kk8Fq�Jq>�d�I��h���t3GW���>��8�����8��Ktb��Y�n;f9�����&��T�\�pυ�z~v��lv�2�%q���&��nj})nї��ڪ^)�EՇ�H�lh�vR���~�g��%�޷�	v�؂�������>�����KϿ�� A�׮�z5Gܾ�W�uOo=W�'/�\���Y�r��2Z��V�GPy���a \��-tJ���>A&��!�L?�<n��.'���"�ٽ��=ěBs�����f�j`�>�SD�.~t�c�1�<� �Q!�����0���D�o��@�Al�!	,���u�ނ71���CN����̸�+U"iZ,�}Ʋ�2%�����@�RN:I�D�o}�6m"9\����q�-����J5�rDX\��♾�5�I-���]�^�pI*�Ajx%6~�w�G����:[��S��  �C�{��^�N��:z�\��hq�5�-q�+�\J ���`'a䜈RG�LL�\e
��隱�d"��S��G��Q�\���;S�Ly�蹸��L)/Qr��t�H��O���!���i"�ǁm;D��ů`7���R�5k5���y(v_Z|&�3�y��n��\݄��*%z�/���6�oa�&+_���зLr�Y����ۿ7��:?K�!,�[栙:���J�Smb��8�q�)4cˮ�v���~I�_uN�3˄p&� ��ram ׭߈j��˗'L�^d�}�+_�#�=���;�=��i�6�bjV\M9�j��x�<����8*j�
��^��D���	�AQRƵ$3G�DNX5)�\&��S�<���6w&�Q18����i�X�ȅ��G8{�c����]��;�z����>� ��&�P}�Y��X����\<qA8�,��]'Rt�=��� �*B����(]���0����8��;v#ĜUK��!"]91�>��b�=c��f�^��z�ʈ+;J�^���k�sM�	&̑�j��w[��Y��:�� -�O��,!rԈf��ݬLO#�Ɛ��!�AUnVB��)uY[��	���0��u6�Q�cM�ۨ	d.]m4��)�U���	���+ j�Z�������Lł��Ċ��ڴ�5�K�4ѽc	��!� I#�G�IZw�Hu�!«�ذm/�z]�P\�9�N�ئ&p��!Ď܇s��"t�6�68��7	;���+8����@51H��<DQ��㐂<0}�d!����ILb��G�>��^�um6Y��[�1s݄�9	�~]���V(+��2��w~����ы*U���%q�~�q/h��"�q>�f�Ԝ�oI��10�V��èx.�oߊ/<�0��ۋݻv�^sq��G�������3X�f{�I|�O���8���0�(���wU����~o<����г$���`��W{���SȚ�4�g��Ĳ�SsŚvR�� �@)"�H2gk��j���@�v�>vG��]�VD�v탪��B�ew[�v�������?��/�htffP�u<����&|c��V��6s�2�g�Q>�Zp�X	�B�V2"nYu�ɗ���<8�

/�V�-�u�R>�y��NWW�"�x��npy����B��6$�':��!hH����D��-�|��$�ڥ�6lD��y��围��&DDnU�JD�EUjں�R���L9���ښ{]z&%����4f�1�
����R�L�H�����A%��CNV���oeKMF�{Rv*`m��)��3h�7��ʍZ8� 6m�����P
p��C�"�GH��>��g�l3y��u���v�@�6���Z�Iy��۾��8]<jV���Ǭ�ۜmv���l������"�\�d�eK�9���s�2 ����V�:�2����:һ���As߾}��?�o�w�LL4q��A���~;z�?� �v!�ν��>� �;rD,�m�R�*M�Χ.
|#6.1��p%	����B�5�_��Q��)�y<�G�">1���d���Gq��>ֲ����""�!�{8,����Xɒ a�o�A�K�U.���Ʉ�M��X�[2� �?��Ta��t�T�tQ�^�j���ps������H�O���k����"�/k�멹��y���#v�5��H졉,h��h!��V����!���IbJ�k�B�T船�WHD������Ж�H���y3��Ţ�b����vɭ0�_F��ک��r���~���v���,d%�"C��Գ帵Teƅ�:������A�%��VB��!b�1���/M8&;8��hM��.`+�Hŉ���Vo"��X}S�alkw��ً'�&,}�"���L�+�"��X��6F!�sKJ6�V�yu݊6�>���g�	wk�lqX�̡�_J�fYNF략D���}����^���:��o�.�q?��Oq��{8��{���D�:����*f�[��֛����a���Z���M��Lh8>�)�:�¼@��MP1{\��f�B4D=�9����S�n�ND��].f+� �¢�_<��_� �£W���B�底�uw����T�8��M�\S3�����hL�D��epq������z���P�� �:~g
���ה�2�]��UB�Tq5����yƴ���'q�+���ϥWʍ���H�f�41��>\#�̂����7��c���u����!F��QLu���1x;+�A$�B����zM\�I���O��9"����K����.w
��^�c)�erN9-A�o_[��RJB�"�z4�H�H�Ѥ�ݽXE�:B�%(�˝]�̉St�f�HrH'�'㗐9w۽p�#e£��<�s^��2UB�B��}���0ʐ8���:o���غ��]�E�
7`h��aI�2G�f�V�e" J�]����eP�Bʩ��fq�HYc�+ϳ�s�=�����Ki���B�֐O��5����T�LNC��\�kl��[��Rq�)f�����?@t��8'f�X�|-5�S"l��&Z�$Н�p��dwZJ�,��O�DA�?�̑�ptr�\������z���+v$\~���}+V��?���)�DbkD"�\7&r��HL��cܦlccW}l%�g�
,����͈�!`�3�T��s��M�3�!�'�e�������+�%׮g݃��-(�Y�i�C�w�������TI䈵��O~����l��jT��������W	&�M"��Ūǟ����Ȏ�rV>��\b�R'\�5ws�2)��]΍��-
u8����Ij��!���9E,�	̚��B���=p?-�:T���֛o�}劐a��x�.^L$�&+��;�-�3:(�6e��#b7�i+Z������Ӣ��L�7Ѹq�>���>�na=���YȌ\��]��ú�x���
�e{ӗ9�
��2*K>5��b�����hZ���1�Fرc����[M���122�f�-V�N��+����ڠx�~*ǟ9s�qz�%15�g�2S�Z��G��{�Z��g�`�p8���`J����t���%63�@^�5%!V�T�3��8���10���/=w�n�}NX��.ً;��x���4�ܭ��Ћ�$k�1�#&t��u�q��;��zn�)�|�؟"��]��Y�T�!3Y7>�eAL�)����~7�*�N��sll�y7ñ\.c���u��5���3Kޮ���t�w�΍�$�����O���a�#O`�WYYd���9����8��aIq��}��{^l��T*h�y7����!����z���PPmܖL0Y0g"�=N��L�ܼ�>�IH��p@=3�I�dl��j�R�\ϖ��SG48�V���օ<�rp�6=�^� �F[��ؓ�	�(�t�
�`s������M�^ZȺV��n�է��]1-�'�b����e�U��!M˰V���I���K~;���jـ�I��࣏>O=�������sg�˷ߒ�>� �4��[5I��e W*$$&#�o�pt/Y���$Y!7�i������e�pp�{�Ĳ��6V#�¤���4���2g��/��D�輧[D�#4`�.���˯"�߬l��W�!�Q��r��I=�F��G��W1�ĀKgh_7A�C��d�	1��^t^{	���T���$�9q<����F�D�2F;������3!�=b�nSG��zYK�{Y�ɻ� s�1j��U�����aW� q��I��
ˏ�l1����h��).~p禚Dhr���!�n��u�[�A�b��݁vhG�I,5x9{�Nfdp���f�R�8���Ҫ�a��KRE9O7u� �|A�E�iv�jDĘb"n����A��#�x�(Ii�'<�����c3oԉtf�%Q�xL��!�	�Ӝ�@;���s*k�">y#5qn�G���Y����6�7�J"��?e=O�3'{� rw�(���Xv�$nكkHrOW��vu���7��fI��6�ܵ(L٥��	{��¿���
���l\��uy����w�����A1��U�7��f�<�ʸ��"��t��L#�7c�.rO#I;^)i�)*��b��$��^�:�X�|��P��N[4=C�5:׏�Ct�Il���F�����q��T���o|��S�4�\!�عD$��%"���G2*iy����V#kyc���mܿB�$yr#�"�$�2埌��\�UA�#?BK?/�pL(=�:�L�=�P���n}Q�I$��$W�$�UIQD8�,+"�I�J�KL�3�2!A�ct~�Ϟ���ޛ�u�gb�Y��^�� ��"EQ\$R�.˖=�g�v�?�I\�*WR���jR�T2��L9c�$NƞG�5�G�D�I�w $H ������-g�����;�\�mxӧ�O������{��gq���A��NUȳ5�@k�:L;���֒/����J�@���(<Ny����2����'A��Ա20(ѥ\gM�C2>t�f�wk�F��&h�~�ۙ�#p�� ����F*��"��&=�|n#��z�D9��ԑ�[� lp��gϝG��)5x�E�_��ڧQ-W=��e��cXH��B�˸���KQڜ���݀e����ˣ�c�X��y��v�A%�Mw�EI���^�~��ugN��~e�2q�&���h�Z�lq�����Y���[��*�3�ӹ#/o;��E����1>׬���?%@�L"G��賀�V�ϕ��dƍ�R�)(���_�Y!B����u�Q�=�����9���~�� ՊD�r��n w�V�Z.�wۋh6����@4~�������wp�"qq�7~����U�f����.<z`C��`6)r��X�YWϓ�1��yE�z�tD���d`6���ř�r�%���R�Jo[��|�U��Zs>��m4�z�6���yS?�f�'~���Uq��4c��Ԯ��� 䑰�s���>���P�D������ZíaL��A�=⢊��c��.�n��j��Wю���tW��Y]E؍��,_�.�����#�ޝ���-�֕�bj���v�۰�1m2RG�R�,���3K�0���9���I^��%����'�����o����\��Sze1��@ ���69(�L^���E�� �;�z6%0�(�tp�8B�� Or�hnP�A��\,W�VV@�^<7N�����2�xQ<�'�����庌�ZR�D��駟����S{ifB�޳,��
�	-gΌI�q~Mf�\ߓ��-� |H�#6`j/�4��J G�)��V���I�S:jṠ�+Z��Gϭ!!���4�����������8VC'�O�F�-q�?����Ѓ��۠Gd��Ȑ�b���hO�� #�^�@���oa�m��ݨ���)�&���Ʈ�~�/<�^��9Y�a[��`̞��bs��UW�fuh�V!Pn��V���^��s8�hONc��$���I(�,�*wu@ �k�f�=��Y>����2��P�m��o|ހ�|���D��Y,���G�Ve�d�=���f֢(FF@��:l���Ċ�Gv����z���,������mh�Ո'�.j�\4���j4֮�ۢz�t�ZS |�Ô�Mb�������	��t��0�}�=�aL����O��׌+���<
#j�9�d�k/���y�y�13:�kvߌ�W_F��Y���4���\.q�G��i�<�VI�~�cdLB67���S:؃������~�.�8V�WV@�^\G�U?�����1��ϥ�l�o���r�f�k�,��Y^D�V��g�����X58�];w`��M8E��o���C�9T	Lp��r��0X����y]]
k�(M�C����|O %Ord	�IZ�=���^"��f���,��\1�9S�mW[H�A��`������8c�,f����Y�н���ǽ]Z;]t�.B��Z�}����A`�u�6�ҽ���<�֝o�62*��MqQ�������a���#��@#�`�s��/3)i�YGfR��	��~�$@T@���X���;��9�6j�.���Gg~�TgR`������b�$-�C�B�:�B�D��jeS'%�t�'3K[��z��:?���q	�Wo���Y(V�}�^'���܌�_��I��D):�@�@\ڣ{�����wG�������^�YA��D����f��Sq[�&�*�)��@�pnj$��v5�C�V�Ǫ�vѭ����q�#�H?�t�1uJ�J͒��VL���	oIm�f^�۰k�Y����Q��:Mz~�B�J�v��[?��7
���x<aid ��l���,�l+	�ia��Ǜ��>�̰_O�Q�����T>�N��F[� �*�	�.��4,����xA5Ւ��cZ
F��]����1�9^ɓ��]��)bY��%�4�q.T�e�����Q-���%O޻�Y��|SDo2�K�k�^�c��x�f�j�3z�dx쥓�N�m�N*)�<Y*�B}&�I����h9�3��!��-�Ш`��-�ڗ���~����_���W���sx��q���Am�B�cVF��]�+�K1劫�oƀN���j=� %�.�"�}�j�4eMs���4�	�U���[��K�l�D�8���a�׾��~;�Գ�g���K�f��ct�.4V�h�V'\��`{�8��
-�Q�(�9ss^Gm�`�"lZ�S�ui1Y��g�.j��7�w�N�����, �V�00t�d1�ڢ�m݅�ߏ�������[�`�
$l��HgY�+��{J���l���k��y�*&0�Cwr5�@�k ׇF����c�>xHk�Q�3{�H�c?�-[��1�ë�!Zw*���/�0?1���A���k�� 6J�W�,�b�#c� ���#8bx^��Nm�ej��f|�V$���}�m~���s�,�T�X�� �ڵ���T�Y��G���q<�iJ�V��-I�*��u~U�����w�4W�C����k-`�T7mFt�0<�`x�2e�L
(�L.j�3�ttj_��(B�Ƌ��YYG�ah_�L�v�v	��V_V���+�K�z��W��eqS��KgO|�O�,
�<osvF�;���E���;:�ʕc!@r�v�H^|�z/9��Œ���z����K�{)-�L�\"��.Jj�s8¶�J�]�Y��:ʒb���V�o٢��`t|:�E4]-����������K;���,*��Y�����TJ�-��Zw��#����|d �	q�(���o��_x'N�c�@�@��M������|���3LL̠B+;w{�=f�K0�
���g�1�ʭw�:4�޳����8)<�/��Iwa���у�Ϗ!�E�c~��ඈ�T�h'ڸۿ�U��AL`�:����-���O!d	�7�Ӧ���sa�eJ���YY-��z j�8� Q��R:��0���b���1{� �9�����6��X|]}^��ƚAx���q�[9}T�r���u�o��/<�3s�b�L6�23����� �d�z�S���0�,Z^��G�q�^��!��2U��q�l�M��<��,�:�dfA��k�Pٰß��|��pS�Y|Y���,zǏ �ܲ�I@n��a�u;]�%i�f��.���q��:�=�S���&�"&l5������>`�.I��C��5�G��%,���`	�w��W����=�([KW��R�>o�ݷ���T{mDɼ��4'���Etqt3˞�0�	X��>���9�u�X䌮Yrd�(�7߄���xu$�~��)�rQ����D��+���˦�ޢ�E��T��\1�+��/{��!���߽�����םe�'?����ӧם:ujk��&��Ѹv�$	���n���T̪3Y���~N��Se�Ş���5Ƿn�������UX.{����mN��'�^{�S�6Y0#��-�Ǡ�Kd[�q��.G�N	W�MGN+wx�;�:Cm[4���au�ؤdؕeXMG�)��]���dص�m��x衇p���7��'~�?���9f�⸇;n��}�x�?3����4}�m�q��@���n=��K&\X�����Tw'��1���8����SX=v�mү��-,�]47���/�`�Mw�{vB$-j��c+]���'��쟤z�m�d��(SI ��I�E�͙'O��SOc��u�����	�`�����݄U�6aս ��(\D��(&O�BtdذX��f����n�J�$>�up5W��;%Y�m8�%�s�I��+Lg~`)�D��s�������"���9K��z�!�6oE��[h�s^82��7��{��I�U���6�i���N�{�]�������ǥ�<��<����׳�}��vj���v"�v_�1�}'\o�$��ql֮#G1O��i��(ϐP��6o6m�;9�?&,��8�ɣh�Àbaf�oΏ�S�(�z�)��cd�i��da 0���Ĕ  �u�t��)��i��
]��]|�u��m��صk��f?L��8���Bg��1v�<�:�c����^�#�j�Ν[�رѷ�zk�ɓ'?�g�g����n` G�٢yU&6*A�^��沀��;t�34��+z��*,��D�'Y6\�YExk��k��t���ѹ�������|$P��	Nυ�;.{fw�ю���;(9�$��u)-���}��&:�Ech��~�eIxυ۶=��}{_��z�w�����e\��*-��	�K\�B��@�6��0*�/	؅��u��f����vV���NO����e�mp�R�g��\5
O�$(��߻��2m�t�2m(�^!�w~'^x	>�f�ҿ��*��^�A��8�xx���na��w���,Ji�45��*����E2D(��5��T���#P�zݵp���s$g�Cu橯"t%�����T�
s-��es��\� %@��Xgf
髯�_��Fy����YЛn!@{��\����ɪ�%��eE�4���Ϡ��c�$&�~�^��9߻�F��ٶ��]U�**�I_�#��n|�844֫æz_����}nS?y��~D���_���74�af��q�1ۘrc�	�l�����	jt��AW��_�G��D���YÏ���mԠ�|����O��Jd��F�m[1�a#r�/Ρ˽�J��\4�
?8u�+oG���C�����o��T`�bO�L����"N�9������|o�y�n�j����C h~́�#G��8qb�[��/�⾷�~��SSS�	�fY6D_a�M����-®�����е�t�]�ϰ}Wݪw�A�Ji��i�*O���?�w�0�K�P�?�Q�v���v���嶯R�4�<s��;e���5�hgaw�?K�_L`�<��b�.��e��׼���56����j�V̸u�m��/�����B'J�2k�Ѧ���ʗ��2:c�@�S��9)Un�g�	-BL�R�fK���|�[J��Pa��A3%��Yc���h�'Y�u'_�g�6�lh@��\���v�ŋ�e9$�ft���E�ϢK e Հ��켠��Qa��@/Mp��ć���O��`lLwWm
�Y��9`���z���LV�V��"��m�ו������p��1{`/�yTR��҉�S�3T� �<8I��� ��T�F����ۆ� ��Z�~p�t}�K�dV��WK��݌��=3hNg^~sϽ�F'�9��d)�-Rg������X�~���e�e��,�7����4�:n�n�yg+�������"N��V��
�'竍*UT֬���-�����S{/b�%P��$�4Z��M�#}V��-�4>��p�9�x��±'��st�A8aE��
���uھ��:NC�'�*2ԕ%��O������F׍;]��x�#Ouvk��1�~���s��q���ַ��g�{��l]s�gY�����:�Q\e��_�����k���Z�1$VA�GG��*��l*���ؐ��:�Ձu�X&�J5�Qdth�2�����E����"Z���,�WW�� ��'��/�:FKV���ٙ;Js�v[9~أ6���8*I�ͯ�G��^6��'V�*5�����.?�ű�dn��S�+�:zm�q���`ڈ����͠���MɎр;~�8S<�������Y4�lٲ�h���Ϟ��\����lТ��`���	����6p;"{az�榕/E�3_؊�]6�Hӕ�&Z�b*d����g8*-�����ђ�>t>ڙf�X�6�S�9�^|�z#�~]��6,z�FNՓ,
��tAk�MLbꙟ�����.٩<K5 a��\q��E_%P5��e���a��I4?�	�t�u�%	�87��p���ȌfEJ��%�����g0��+e/ғ���-��qV�\�%Q`ptl�h��E��D9�]@�BoR8������Y$v�G?��j��yD�g�7W�6wEj�kIn��5��v�37?������>��Ю	u��h�1��F�E�����#"ׁ��<E�E&O��QZ��M�������y,��y�|�	T��H�p�vhLukX�c7�a�4DDq�;���Ǳ&��cH)k��� s-i6i6�Bw2���ǟx�~o}��S�Bk��v'ξ��3�t��N�ΰ��%o��{�E�ť��l:������B����|1��g�߳������1�*m��Q�m��Օ^өE9@G,%��n����Y�~/�?��x\3�3��t�Ζ��q�&�M]/T������L���
?�Z���נ�ÃrL��w��7?���/���A�\��-4n�A@ �Q�J�@I䜖�x��`
�)�.UQ���{�-��uղ��%I%�Ӑ&��h��S-��X�#�²R.Ka�A��I/CM	<�����XG��`z�8q�W�#[2���$i���^_��' ���y��ي�E�5��	���|SRo�q��b�a��=�ނ;o�7ݴO��/�"��i���0k�y�',�N�%�h�Ey��z�	2�7>!��{�a��4}�T�g���/��a6̐����)�b����4gC�g��P1���1��mn��4��&aĘ����5�>O�R�t��G1��s8�����1p	�{�]�H����(�bVkR;�P������7���;ܺX��@F�@����^���ΞL��gNb��L:$,`~~���&O����toᚦ��{�w���m�&z����V�Fwa����Oa��¹iDiC6:�JUI%��Ӓ(����A��߇1hS����R���C�?��U���a��Q�b�s�X{?������E�V�:p%��>�܇,2N�����/��;C�f&`=���j	r]�N�.� 2-J	��O��ꑤ��
�<��I�,�΍?�f��{�pvغ�vlT�s��c�N�>;n6,y�\"7�Y�7N���D�)�z/����y�!ܶ�&��Y��x;=�=�i���w�y�_�7��'�u����(���t������$�Di0G�v��� Gc��k�Ȕm�����ҿR��x��#��&E������:�<��H�z����_J9�k��ޏ	��E�R� �'�|��eqq�ϝ�(+ݤ�3� =���
������9,=]|��w�D��W�,��"��Oؔ�Xa �n�U�5��wZ|��a1]q*zp9�h��l�q��A��_���~{�얙���C��^|�M|�����ӧ%��0�T�WC�>@-r1+��R����H��p���eq���ƞ	��c�_4g��\'5��uh�D���v�g�!�?��%�?z�@�,bQ�C�W������&�s���Νر�#FG�?�tj8O@���X8us��Ý�E�w�b�M%3��eFoЎU�1`P��������7���qԞy�5k1�m;��[��U:]U�H^p���I��0;O �	�͏�A�ϣʠ�J�u��q4� �MԆK�5`0͌�B?��.��P���欌S�u",��o�ЎmT�m�ͻ%c!&��%`=~��X8s�R���h,P����H�{�؁+ɴٝY�� ��Ә�Y@|�$[6c��[u ��a��6��#�J�� ��}��?��¤ �����0�i��D��=��`x4���/~���/�F�N6
aA�P;/��&z������8�-�4�.v�>~ռ�O��lZ��S�p��G�I�ifqb�G�im�����'������E'�>�����i�u*��3�a�ֵ="\&����������yvds��ho�]$�����V���s��g;�8L�JP�+ʉ!6�`�1�H}�	ib	�k��$�X2����K�%�9^>6 �բ�� nd͞��ԟ�@�����2OO�"��>�b�[�?�pf�4-�
=ڼ�*u8��z�#qjv
�뭟��"����������<�L\�`a~��þ}��_��S��۰��fs {_xo>����F�;���	�L��_4�0�`e|����	�-#�!��X�Ę;�&�����I�&��W�
��aܗ�|�>X�+_c���E��"�)¬q["���\�N���q�# 2I@�=:#{79�d�l`Z����6���Ř��I�d����'�r�%Q���N��sPCB�����<���4��ZU�G�a�k�p�� )�8��� �
��*�a$�K�TI#��u48s�^x��)�#��cs�;�n7GgI���]�ݣ�%��H�����ޏ.�c�;�b�l����#�/." �ܤ��]m�ga��nY�tė2Kz�7XP����,zo�������+/��!��XJ�U���\�Fe���r�D���gدP{�&$�u���z� �̑\����YX8[C�Ƅ�����0��Y�yC-�������\�_,�1M�s&�~��b ��8�@^��MCYr磗vw^��
��p��L�ӡ�951��V��ݻ���*=ע�[j��,�
{�D�7Msٸ~�]���g�H����\���/TU �G-z��޺ּ ��޲5gC�P��y��y��fLE��"����m�r���G}��t�� �����N=�������C�C*�b_��/�n���Dy��{�A΃t���	^|�� �� \]G��!���dJd_1Y� s]���*���̰G��M�Y��H$���H�����ȭ�w�N~fj����x����o3������0�!�*�2	��ޯ�� ��^�:�Q���d䰏R�y7ЭxR$���U�~��-���87��fY�	���SXիb^�Y�� E��Nn�-:�H�1Ny�b���j��*��y$~o��Z,�]qL����>P�ı`���Ċ6mZ�C-�ѵ�	����]�1��R����
0�W4xeڌ�� �#'���À86<��"�:��1\'G�p���yŀ'�����g#���%��x���*��%���1�$�Q=�4����FT�'r�ڔ.�m�k����U��DҮ�ͪ�5i%�%܆!]�łʋ]a�Y9��3�ΰ�]{!mHj�e�!~u�0��>/�b�r�/�<PzQJ��%���#���u}�
:՚��s�M�vB&9�\%%�q�k�T|�ӧΜ֌�sm�S�hP�u�ʻ���fa�)G�Ȏ�p��q+�?���- 4T�_�],x��?���hZ��F�<�����9o��b�q�yS�'nL��n���e�&��ӎ������iy�D��\��q�A�l�&�-ƴsrO�E2�վT�2����볏*�8�b7�Ƀ[�d�(,�/��O&�OZ�o��f����������h�q[���
���1�
�U�sTk�Q�P;M�
A_�Qkf�rNn���D�f�`)Z�ꘔͬ���i.B���ͱ\	0.OL��V� �u5�V���S�v8GfH/5ȩyJ �+�RO��gz)�I�v�SQ�nu)���D�H��=}�qʰ�dV
C:G*����\I��q6�h�hfk ��A�S��+�9ZY�-oFJ�8�`�xH\�?g��33mlNUJR�1�eP��gU�,C�����{���7p�/X��D�h	�'��U��c�-I�j�7�[�"v	خ
uVI��צ2a N��@25(1�;t�(�Y	$c�/e�im�$�q،�fu��,�f|^��� �Ռ@�O��&3EsHιn�P8�Yj���#���/=���awu��^{1��^�������_�߰����4^�����U��>%/6(�}��jѨ:߰'}�_��'-�k=^?��n�	�k��2��K%؊#���f���7���ؽA�Z4�"Ŗ/%w!�#װ��	`�����z�B���
�l�q����ƱC��])�|ئS���&�t�@AqA�"f�-�M�U���ެjى�\�,*�"�aUظNw�N~�H������<t��[�)|���|�3�Hqf���V86>�������x���`��i˜q�(3X�΃���uq�/�d�,M�J��<!��(�8
�`���I(��f������@�D}e1��:�	�+��̾S9{t��dRc�7f�\���af�#�~h�N���0{~���.a�3�$��V]2)�<�,!|^�+1s)N(� �!6+��X�T6��'���)ߛxh�L"�k��Sе��S�l���ŏY1��-�;��jp	�w�D�PAݓk������l� M�dy����5Ix����%���<�
����i:1*�	�vϭ�\^<�C;�����Hhf��\�*Ivp�S��{t��G���pë
�Q�	S4{�~�#Q��i�FbZS������]�gΘ��מrU���ʵ�;F.�-%�J��c�6s_���еi�/�W���V|�+��[n݅F��m[6ȷ�(�b'�?������/�8t�_�k��N�q�Z�*�Jɀ��,��f�$����R�1e���C��8�UtD�١%�r��
#.@��>����qT���\
�8[.4�-Ȥc|5j�q��:q��D��<��7�wJFҥg�>'+�QV��ƬD�-�hǦ��;=84�vR�	���D��bMO��]���+�JM^�8��V�E�����4ڴ���ZV�Q�J�^�zE��wu���\���h�4����V��i�{\��`A�|F�c���)�b�-�I ;e�)-��{�ne4��*���
�`��f96�&)�@����XY�<
x�v�A��eW���L�'@E��b-dH�fK��$���o>wUI7����Uq�M��C�_�>16g~g�	�QA�$:u���J �#��IX�[D��)]k>�@�3̑g�\-����T���T���13�:pH�|�L��8ɵ���1�*u��<4fsy�������_?kl�d��'�Y:����q���[/��AsM"]�D��,�,��"@@c7�`,�¾q�d�P(��e�fM���\t	����������ǏܟuD�԰��~��EH��z���y�#����?�Z�í�쒯ũ��������?|��]�6�饱�^���*
%���1)��V�Ǫkm��v��N�+z���x��̈́��36N"�]P�ϻ�3�p���A^�h7��F1��-Kͦˋ�L5��U;R.+���O�$e֍ 'p�|�l�� lR��~nrK��/�Ѧ���Q/�4�ǉ�#x8�'j�<����T��^��$O,)'��xΟ?����������|鋟Ǘ��E��/����G��ǽD9@��`���<�,���͘���&:�]5/�l���2�$��,=�J��H����|�hP��G����E�I;����f��e��<Փ�/)�8�� x�;�(�jK�����M��]&� 7!qb��E�Q��џpC��cpǦQ2�[�׳�\˜߀-�W-V6α��}� ���V�3W�=5_ur�n��\ÌA�Pn#��ns�� �f��o��)����6�O�2�{�6l�.���r��$��
��a�f�rMd��#~g�G�0g��ז->?���It0��)��Q��5ÒanQ��Fl�y�L���5T8�BK�8�r���#�O՟w��� ��a�����ӥ;80Fi��������o��{xy�y���u{:����B~���v�'�=��bV:�$m{a͑�!�>����6�����h&*��G(b.U����B	p�~h�^�̫�!l^:�.�i�T��B���3�_����9��4�_��{������)=�X'CN����HH�.��
���A+�}Ի�xT�c$��h;�)+�YJ!�h2�����f| �h�k[�Wa�X~� ,����R�$�p��118ԫ!x[6n���$N�8���)z�!��<)q`C,�/�\��u��ׇk�mWk��-��vF��h�tQ�F�L��&Z�o�)�Rgp�	O᱐�r�T/]�,�2�d�s����,��P��gZ�Z�?�o���^��M]�~�h�_m��-iֿn��\���LcJ��=��ߥ���_4!�)��|�-�,�}Xܱn[������EZ�M�^����Mf��0C�%�ܿ+b-�qLwL���vw�㪸�軦}?z�)�F|��hr{���rM�@N `7��'K�x*���p������8Ǣ��ë�jT8�y�>#�7�}���kk�	��+�҈���ȵ��7��[�C���eR٘�໓���S��u���~��L�YB�#��Ŗ��;���,D`�׎�Yv���E�Ck��,d$��R���A6TYV��h�\}R�ı��'^j����=T��C������ݣ6{]���-^sS��Gh-<�i��SU+&%f*�9��Ūa�,_|�k�1���wߌ�bժlݼ�&T����������^D행i��vDq��L���|�����9�_��*`I��BX��df�c�F~p�a_H�����K��e��>�AT?g�꟠�K�pJ��L��f�򟾭;�o�c���$�ka���]|�[��GBW�)��_����-`*�N�Ӈ��x�V=e�7�F��sQ�V��� ͣ�N^� ��F�[a�ڤo����#� �G��l{�7z�-N���ҬE�ݕaZ��y�΋��}'�uql>���!��$��.^�{@�kM�,`tt���<��ؼi=���]������(N�����H��&͓5#_�L������\*���h��)��>�D�%/�?<�1�b�q��3|�#?�nE��g��
�5t;����h�&Z+���x�@��%]
p�@��Z�G\&�[x�:$I>�������rٙ����*a����r�h�9T]�z������3_9~ȣ6i~��w}�(�T�*N��r��1�ݝ���@����Q��um�RE�����@v��W��W��5|��{D���h�imϞ=شi�$�X~�N�ufzK�����Jzѝc�8�=.�m��!�$���"f�ү�<3̘+~k�4�A�c��Z�������M�Y��*�dQ����^µ�v͂�A���-�ɗ�D��E��,��99�lAJ3&�	80 �)��-`�d}���ֻ���*�a*� 1/�y( �* ܲ��`�ߎ>KV<��Z�����\��Gж��"#a�� k1s{��5�2�}M2$\��e6������e��tJ�"����G����U :ǥ��M�G�����ǎ���^���G��ǜ�B���nޅ�[6��Ԍ>[	�M�ռG��J���J��)��*K�*�\q�p]���y����d���L��X�U�G�7���4@�ܔq�GN'�B-p�d�V]�\�Mt���x�ͩ�w-��4�j���fG|jԯ�֓8Ҋ���#��Y�]ܶ���R��@J�$*�>Oi6?�E���\�
�g�/?d:A�5��'�� ȉ�s����tF�^���6��gķ��٬ȃ>??�nO�I��9ubj���Z��##yA�� c�e�,��"���@����}��!/ �d0�Z>a�f���4 t��@n�F����n��ϔ��)2>�e�K����=j&MgL�����q��(Ui\){_�ԯ�μ�3ZXP�t����Y���q���&�2[���� $���:]�r��m�~��K �#.�˥ ����2�t�1$=Qp�u�*@`8[ �QK^:��M+��T����Rv�`mC1�BG#�"G�s�����:�h{_�/�Q!�U���qaVe4�0�\���A���U!W�i�ۘ)��A)ɪ����2$��W�i�����Ly^�Hs.p,�әU&�d��jh{�N�T�c��K��N�̦��C`͉:=�m+�V/kF�^�Bc�*�K��K�����Z������ �7�m~��6�;�r$;� T���J[$�ۣ�&.���r�uU��v�4�c�[�
������J�n���:iRVb\u�9�Ո"�a�œ9G��L��'�?��}F��>�أ�o��7񳧞��ܢ, ��1�86�N���$ΎN�ŋl�>OX�%{f#��;z��ͬ���Y@R��\� G��5�� ����MJ�e鱖
{��Y
�Pf����2iKϡL=\��%A3nT���5U[�X��lH,�,�&��t������|_��bU�,j;��d�h�LS^:1L�z���I�QV���wد�5���������7Y�}6�q��M�6��=���dL��ed��.io��,�[�q�8��:)�*Z�R�|!ѱQ�C�H�<�%��)5 �]�k��S��.7yd/%�s9�~n�3�ukY�9Ym}��u=��S���̉UO��� ��n��+�<��a¾�0�g��c����	?�E�_l6^���K��q�` Y�>���?�����d�Y�ԋ:��������t=��^��M`	c�S湘��+Y,���R��nL׬z�w��H� eQ4��A�x�j��_9^��k'��Q�ZE?��C����z��K<(֤��Q"g����.��2Wf7��������i!LŜ������c�=/j���Ƣ�������W� ��v>�8���>�w�u�碜�X������Ƃ%Y���T�O{��YB�l6,L
��%���E^X�`�x^���c}���%4�fBx8X��7!:Ɨ�|M��Yd_�`�ʦRU�k�d��~܂��׷M����0�B��ْ���˳�$1�i/O���y��7/��23j7D���e�d�7=����l�!�d{�����,l�"l��b�[.
Zc޴@�1 �h���7���dZa��4�UX��'�7o݈/��Z5L�җyq~����iM.�4y�t&�EG�z�ZK�h�Ռ�=qZ��۲��WY�g�쟞^�&�oV��YwC'���q����k�qoM���H�m�*�9�%A��{�������0oL����~C�ϐ���S$ ��]�1���eV����ш����(ӊ�^�����q�	���f@.�A��~h����C��D'�v�{q�U����J{n��}�Q��U=�b���V�3S�я��i�#�$�ެaՔ[��R_&=q�Mc9�M��o
tQD{��ꨥ���&Z�}(��)ٞ��ּg���T�1a�/�Q�����!e�g�`-9"���({�����IS�GK0b�ǂ���2/X.͸9���l�Vn)z��.}`�ϛ���i��B�{8��m{�\�ri�r���_J��5���4���UE���N�%m�*������V�>��w����;��S	����]�XR�o
[�����)X�����g��|J�+���
�E�[v��w��V�Z�U��u�hцU�4��+w���l����zv�y? q5ސ��E�h>�k�˿�w�:I�����h�W_}���k��q�o��������6��[<�бz9��n���L�x�M7}4-��\.;�cEm�
�>'؎$�K88A @�U���/+��%����?�_�91-�&ևc��e�iE�L|���ak,{sm�/}Y�e|�֊��]�����w��Ok֭ŝwމ�����`�Bj0j�s����/��͊O@p��H稈�.� An�"}U�ڏH`�)�p.�%���qtj��,��Nf�̇��AY	��c~S8� �W��.Jf]]�܀B�e�>;#f~�f����S�,��ǖ�]O�����(�8����t4�l������D���g|L��O\��#bŎf�G�Z�!3k�A߀V��G��%T��<�&�(YG�o�U�;븉Y=1}�����:�ߙ��n
�x� I��P�u5 ��h�=�����#LE�.s4XK5[+�2�4v5�
2�0��S�Ye�a2��(�C�Žm�~M!��<;.��nG}��6]ܦP(�5��^La�&��aˆ�X�vu��P�Ԅ�c\��?��>������1��i�<I��kzK���Y�n\�d��-��l�]�sZ�����h����Ϩ�ڻw�������=L@z;���ԏ#���YF#�u������+�����Բ�٣[:��Ou��u�P=�p��w�� 岃�JX�g{}�v=^��YT�,C��,*�}f`�xَ��С��}�C��,�W�Kh.�|���!���l�c���:�k��b�ek�.�������8�/�}�<�0���������SO�X��׿��;����8������]`~qN�+|�]Ur�w�ա((-�,#�_Y@��+�Yk��O���稲3}��}�td�ɢ��SFX:X �����4H�/K�/�&"ш��Q��ngar��=P2�����P�$���p��`P���Rm�4 S�@��"u�FI��vbв$���(0m��K�������4;��3d3D��u!�)��N�|�z쨞B��*Mϥ�I���`۽�X�E��]�<S��q��a{T��.��KK��qR~��G�S�����*���g���>�f�}�jnE ��`�L�XB��5��>�k�H�+�ǁ�\���r��{l���-��������^�p���5����<����q�*<s�\���wl��<��U�����3mP�A������|N�h�o�X߹s�/q�����4ܟ���'q����;�Jh��䡒�_��\�$ʡ0<�]C�x���1�{�ZRԅ�i��· =�C��\�|��~_~��~���Ӕ��%�'Q�4}�SJN��ӳ�"��<r\����L�Z��A��v:[۝HN�Jv�Պ_����Nޗ� r���>Vf��E�,����_����ǎK����'���شi6l؀3㳴���C�s�&%�%罔�P�;�^~M��bÀfu\���4����g�\a����JU��؏:��2�?�x0�Pzs��,�rO�D���svn��iMQ�ذ�%&d�O�f�cf��yO�Q厩�#�9|H����#u��|o|��6��qRX����6��m6�՚qS��< 9��<�>���]�0}k��>m��9��ag���B0�V�d���F�t�a3�3�,rw����Z��K���y	3f�A�?t[�1r��(h,tK�Y��1p]k�Dl�o%e��p+o;�����?����\a��KU���z���G�G��p�J��{����r�A��M���/���Ek	ą��#��:G�d���w�E�5BX�ec2�:�k�=}Tt��)ϣi��5���M������2�|��Rl͇>��k�k�.]/ϝ�x1�����=����Q��CNQo����l�j��:�R�}`ί_���^�<R7�=����K�s[''~�ĘA�U�ɹts�x���jkP���\�����`o���#*M�}�vl�4��~��8z����dV:��y���o�:>u�x����՛���Gs�a@��S��8�ی^8����m���x' ����xJ�izQ7���k�٭�WD�j!c1Y�fP���P� /�c�R���ȫ�g�9��J��v�ٛM�b�U�=����bJ��1��G���=���-�&�fco����zߙ9dQD��Ln�e9�[��B�`&���C_���>��wv��fT((&��=���~���VZ�ܳ6�K�mKSz��`Q�4j��ozF_��*����U��7�&�����&&���������)��Z�� �����w�[)��\v�[��[�����R����/��_|�׎�'��v���a���z�(�k�{���t���Ր㩵�����12�����b�ctx���-�f+�е��H�X��g�,p*K_\LYn־�)-�V���O��B?'�6��A �5K����\O`����&���s�	h�:���	Z�8�]$��d������lʹ1T|����ɀD������~^�^���2��g}q���}�ߋ�&�oK�����V��h��`���&��-��p��|�0Ӿ|	�O��&� S} Y�'�B�ȍ������h7�#�<6*f!�N���K�,�7�J��P�ִ�����ʹU��4p~q�~r�qpR��m�)�:���/�6f�_�*p�ڱ�+ �,׼}�\\���Xh���ݬ��Y_B�=Z4Tf"�oF��^^�3N���7�''01�����8y�$�~�)�h'�m��{cl|/��W��g�10X�\�W��%e���]���S���_�f�T��������{��%$��RZ�;���\�
���)X�\�>ۦ�:8��;�hY�V��ѬE ��p~����i�L���]��
G},p����Sڧ�����K�P�����Tq��ĵ&I]ׂ�l�	�F���n!��$����~ny�df.04&del�e�R����LY�k��wPp�ێ���¾�>���,E�Zp�+u񳎩C��\m1���Yk��+K9����C1Aky��+�++ �/q���:�oI�!�i�N3�!��@w�R�	_���.�(å�������[�n��{�'�o|�7D	~��L�Fx���w�~p�U�Ձs4��"��勯~?�~mE\���8-/|ykv+��962<��q����1-jө�ruu 3>�DUZࢣ)���]���f�,u@�Ȅ%�tdi�j0h}��]t=3W�D1�ڀ	�g�Δ�{�
�Ƞ#`�����F���M;4<e���¼�9f�ȹ���<���և��]"O�(�g�Q�:L$s5�ӌb(��Mp��3YJ�Aͬ���ᾓ�\��[�r�v�OR��E�L��Ɗ�����c��(T���(1�2�4C�u�5�eq��K�Li �2"*�*?p��ɘSť+�++ �/����V��.K��*��7��+�Z�/wݵ]�CRٓ��%�	6Ϝ;w��ַ����ݻwc����Z_��&^y����؋$+��tI�wSN�T(�P�m@`Y�/1�f���� ��3�-4)NV��iH��,`��$��R�u���#�hӬ6"j����m� �v�T0F᭮�� /���j�I�������;s,��A�m�İg�i��;�͆mS��_�0f:Z?keuu*'��h.��jY�^����R�ISF��F����9��6�-M���T���Pq����;Y�+���� ��i�i�ʜz!��70;��=ĥ�)�2�3*�Qq}�mD�R>RYq7x�<O' ����j�����`���v�:��l��#fg+���i#��H�o��:N�<��7b�����ǎ�ԩS\�C��J�R���x�Kf/XXZb]xq�3Y�z�Ne�H.c�_��B�н3p]�A��#�%!d1�<�����L$h<�����,B�o����#�т���
��G���]t]m�d�A�.Bj N[VoT���IW.����XL��.�s9&ES�=ڀT�3���^ؖ$��~����t7@i��>� 2�ʣ�ҍVs�H?&��e�/�Q��
����%�BkE���H���8�	+�*+��Q{�Z{�e����ڥ�>1���<����>cAtI�Gu���r���W�e3Ĩ�Upg	+i�sD��P�b�t�+�Z��r��Y�J`��nխ��j/���M�6-��>���Pƒ�v�
�#����G��ַ��Id���2o�^�-�Z.��.+L�XV@�^���s��Lf��]Lj������$\F� �'{v��\��j���}�j���hTk��-��a�:�۷'����b��*tX���So��M;���K�dK�06J�J���ٛ��)f��JCk���M,2�g�mQ�b��[�F���@��:�gpl'�@�8���Uѡ�2����v�h�ҮmXgm�=Bl��;�e��o)�ӵ	Tdک/Htv�6����*�%��h�30F�y�`!�W�"bY�6<Y��t/��]��zU�_�8����	]$�k'�,5�z�� \�^�KרҹSTk�
���L�a>v�1�@3K��,��V�h%���j>0y\��]��H��Z$6˔~G�%�]�y��0�3�.�e�����ȹ�D[r]��S:��#�3G���;tM���qnfZ�sRo1�j�.c�Ӌ�^+����"�} WT\iT����;�	B)��ׇ?\�(툺Rn���V�usYR����b�6���B\�5X޽�z�c��G�U-b�6lX/ ��D��n��o~۶�A�=~���w�����"i!$ A9���./§\26s���Bk�.a���X���i<"sT�8�l3c-��*-ҋ�X�9����N�A0�pT%'�v+����&B�^M����\�a�x"0D���U�����A�8������%pَI��F�M1�e�CߌC�j�bV*˫B�ZՐSǥXd�CX����uC6I/E'�AL@1���_Y=��-�j:�Z� �[%`Wa�2B��Y=7~w�wG��>X���*�#K#q?��+���a���.:�ۨ"n�X]�P �"���z:3�n��&*f�X�G���~�ʀ̈́t7�0��u]rj�}n���S�&>u I�Pk���Y��{
5q����/��&�(����5�|1�
�N@Q��0Q�u�L����&z�3ѳV<�J��#�4��Tʏ����렰��
���
���K�K9?��n�U�n�Kw���rd۵[l �dGP�4�:3ō�\���K�~�����wb˖-l�����ⳟ�ݯ~��v 'NO���!����7��Z:ڑ�rmޅN�Ċ�!���m�Q۲��$�q���O�07x�F�m��]7���C����OD`!]��7��('GF<?�l���#G�L�aU����Km8�yf����ܹ��E�#:�H�=��I�fou:w���*�� 0�����5lܽ�m��A1��3;r'�B�ͣi*�e���}	�Ti&�H-n�@5C�Us,�9�w���zl#z�߲ޭ�0��a,�=�:��x(:�BܖTt,��@,�s�)�b�*�g��Qi��GFF���aa|F��e��uc��P��)O����͎���:Xw���?���^��f�g�xt��ʀ7mӵ=�z�Yj�E�����A�����c�h�ȝ�拃&T
/$��F{1"���������
��$�A,by\�v�����i���1�>�e��^\O���Q���TV@�^�<Ϝ�^ʇ��մj|��{�oe�5���<1�qE6�q4��?�j���/�$�.��~4�>~��O����E���w܆m[6c�Λı�}�/]��T$�=
h�$'�)%B��TL�fGW�K�RE}�M�#��J ��L�N�������ç�N��B��=L�>)~Z�M;�����`h ���}l;}
�?yS�'`�V,�_�=�=�)/��[GTVQ�����S�±�F�MPa?/���V1��[�;>� ܻo�j&��5�c�|�5��cO|jq���E%l�B������X��#�c��>yy�#��P]m��& ˦�fo�:�����b���bb���uW|ɂj�3�,&)��3�E?����q?Ɩ[���v!y�e�S�Tc�g�-�6m@�_�=�Yg��J"�t����>lي��#8t�-4�]A�+Q�98V�� �.,c��>hհ�V�� ����� �� +O�l�vބ�XH"8�~�%�4G�+�&轴��l��3N�{��JPh�9�}ϝ�5�
@PYp���. ��\O��Y{VʍVV@�^$���2��'�륈�����ha�hyv=�_�{v��+{������
�3��_���۶m�K/����yt�mLLL`xx��d��Ŀ*����-Y��̆1{�@�j���n	�UCpp`߫�V��;�nq'Nbf��Y�I�!D��]��T9p�u���ccx���^�`ݎ]h}���;;y��ZCk��s�j��ĉ�����"'P��λ0p׭ؼ�}��fE
�͢�#%��ȧ��Ԝ8�C��1Ο;�:��;n��=�r'��ɿG�>H`��6�m*���9@Q�M {��"ݡ�~eP��J��,�	)��Wj8G}��R�$�y�^ �o���8�ku���,�!�#E�j��P�o���� 2�}�B�w6#S������(pѠ�a�fq	���>|P�is�`�.`�ZB����́��_��(E-�P58�͠��N�CMԨ��@�f{��6�i�h\G�Н�`�ڪ�.3�4���������Ϣ�.~(�q ��R�̧"Ms�  u}�G+e�|ز�n�� �P2+$�e�.}��6om�p��F� 6Qacf�ص��,Uk��[�#4�g֢Q�����գزe�0q��0��E+��>��]��.�������[	 �ZoIN��{bNM`�:�q���@۲�z/�a��O�	jM��c�w��%�~j���X�q���p��>}/��{ ����[����;��?|ݓo!����y��oG>K�k�Ju�v�C� ��w g����~���a��;��
G�B�ƫ �@���B�����ݍ�w����é�^�8��i�y�-��X$�2�i*#�1��Ә:t��UX��G	�c�����M����]�h�X��6���&���>��ǰ���5�x�0&^܏��	�NdJ ��֐��]�HЄA`}G$����Uo" z�u�?s[�Q���S�T�tI�Z!&&�bv0�և?��wS��FvjǞ{�H��_�@ �Y�O��71�������܈[x �.j�.m,���_x�'������P{�XC�d����߷0nCt�U;&5��x��+R
?])KE�m�?�ϯ��0���PV@�^�0W�\~/\��x����2Iӓ��l&�Tl��1��!��n��v1�5�u�����������9FF��G�"�>;�;��VK����R>2��-M�ft����R=X0I��	�@�M�/��s���yjuD��a��E�}���)<8�Q��R�z��E8l�'�&��"f;1?�,v?|/��=�ջw�۩#G�x�4F��S�����v0����C~Cت}���������^����X���m��	���i�]�u&������� p���;EI�$�$���t��������8f&�m����G�p���c<�o����m��bI\L����@j�z�]眓���*H��*�=�c���.y�����,�	�p:D��L���֧�B��H��g��كm{v����Ñw�B�P���PB�5���84���:���l ��j��6�@���#����E%�МB��W�7��������]�c�A�g�@udG�{	�ɳJ�K��q�|��^UK�����h�MQݱ�Ծ��	������m6l�̙#(҂����O>,4#�6��V�ٿ����p��a�}���X��N4_}������L�8Bϋ�Uu�ŭ�}{:��K�Q~�>���d0��A�T�������õGmg޸���RY~���`g.�\?�A\.��.3*jf�2���_�2ة��W��P�T�<ZA�&�bme��!CuL��*;�'�&=���)���Za 逜D����3���4���QĲ^lhT�X��d�5N�]t
( h��x�Ѓ��`#�v}�f'P�	���c~�@�_��0�s�9I$��m�
.�N*�.�� ��S�� �b�������ZZSs�D5Dv ���s-�=���sVtMj7�Buh�ע=1�R� l�|�"�΍�$�$n����>'����L�:��wa��=��?��	t�+�y��*^������y�m?v���������?a��X���|�i�|�����e�)�o���w��-`���m��o�ٿ�si�ǿ�%8=���:�2 K�q�B�@^���c�g�te�E����9t��]{��``�n:����,�u����',�nA���Z���/1s�"F�����y�18�c����w����F�o+��{����,|�!p0�ֻ8���`_?�?�J�<�ʉh���p�O�$��G_ce��c^Ap��gBW���1H�T�U|��٧%��<��5뻛�늵�ǰ�=pt�Ͳ���$qk\Ҵ�
���t�bY����Y�ׅ2���d�g��w��]�ϐ�� �J�dy��(WJ��ԡ\eJmG§�w~{�4�|�Ag�#��`�{��XIܞ���B1���W��%ȁ���x����i.�������c�O�I�b&������K|���2W�Ċ@*�6����8����J����V�S��$ R`�
ۥ�s����l{i��r���m� Q��XO���� =#/v�i3�.�E��R6��N(����1w�4��m\|� v޶ �����T�A�&�>}��j�0�"`��h�OR̹(�T�h�1�&�/N �%0���p�^�I`�WP�{am�wcϭwc`�����ѹ
�R7	;ϯL}�2Pj8��Q�Q*��e#*����A��!b޲cFwo��^�����y�t�͠R�p��q��p�p*ex3s��L�
U>�"6#��y�hLLc|�&��V�o���9��1{�<gf	�ৗ��Zd6�s�В�*��ұ	�$G_�7�����e�R�s�p�6�4c7������5(9��eM��� �%�s�-t��yv�t�=��%��.�O�Vl�w>W�RD�n|bu7�w���wJ#��~L�*x��&�Dh1hC@�en��s8���ؚ�������{1u�<�-���Y����Q�
�)�p,+u̥��ގ��sa8;<ԏ�M�q�ڨ&����6�v�`���L��*Mb���,�{u|��[���G<1'�p�*�D�B�9�t�$v8	�T������8 `H�Q��6��U���E`�#5][">-�<�#�t��� �eI�@t�)Ӆ�R��\]0�S(�^ks�/����dV(�oa�)\�^S���2�WF����. �s���@R,����
;&j$�6�R������I�F)��jX*җ����U�\�t�+�|���u��s��2�&�S���c��#"T�N��G�E���Γ�����o�:3��*V/uVw]�7d{��dr�j��������t��䲲$qk\
���n�����8�H�)�s�'ƿI���'�&�kx�lK4yr�#q.���y>�a�$c_��%V�1ӿ��T�����40�G�f�֭:M���L��P��#گ3܏#f�O\_��*U���C�ip�z�c��Z����A���cǱ��*�߁}�<����Gc��� e�ޖ{nGx�$�8�Ո�x���	l95lނ�=��W^�t� dC�a�]����ї_���$F�!F蜍[6b��y�ܲ�8�N#!P( �5d�&]���0el��1���������oE��cZ�N;@x��Ƿ`�]wፅ9�������Cr�-�MLPc�.�L?B��i <pk�r����.b��Y�۾� m?�c'���HO��Fi`��an|��6�ލږ-hM�a��� }��K�	�&���%���u8s�ov�ۋ��	x#%l�e�G����ӐDl���j*�hv����,�5β�To�t�d��z��/-�D�+�>>��P���5(9�[��ѩ˻ޯI�D�.I�X!ŵ�T�5i��%���_2�;5���U����@ K�0?�M��B'@g�T#�������fѣ����������ǰiv����/a��#��8�SVb�}�cd�(�qt�=��P!�Շ����?J�L�pˈp���C8�����W����g����}#_�*F�D�M�>��;��>x��#9p��R���"@W1���ￂuO}#;va��E2��V"�w���[�^}���.p�]���'19y�n�&�g��ބ?W� �6���l4�mI3��#�Ҩ��~�h晐�]�4�E�@f�����{�>8�>�Ϭ��9��s05����!��]� ��hM��&=��B t�(�k�tf�F�c� 6і��:|.��,���`�z��#/6fP9q�g�Şo|	���������%xS�(2@�,�
Q����>�wߋѧ�F�Z���`~��O�:YS�I���bUw��Q��@�&3f-�	�bӺ+�,l[)��~�f!6��Dв�-�`-�"�`�t���kP��E0��ĉ����a�	�5r\2�c��;���I�s[���sqrs��F�9�xb��hK�(�%>k��N�l����ҳ�`���7�jJ�<�.f���y��?��)8�7q�
���t��q~�A�5�al��ƻG�LO#�$�i6��s��o�]���٪T;����<�ʦ�&g#h5�-��?x�^�Mw�Cq�Nlf��6�[h���{�mI�e ;���ŝl�ݻ�6P{���髰��(�5����
�e*>ￇ��q2omޱC�����rs����ph;���@���'1��b��}�dq"0p�/��KG�Cգ�=E�� k�:X���q�/�^�}G2c�#��;����f	 �d�2�9 �t-���3��u��>Em�ҋ�e�9֡���Q�;��L�8��Oc�g����-�Ņs8�S�ޅ��c�z�}�6��g�2gk�������7�Ä�]?���b�Ξ�\�\Ū�&�<��$q�( �F��25�����S31�S ��Y#��ʹ���NOd�u�c��/<l�pes�ǟF�c�1�����e���eER���or&&)>p ��I�?<���P��Q�c�t�����7�'l"��&PR��L�T%eg��Zs�p���6��}��s�g�d}3/>��p6n�@�V;�BcSc�0Hm_� 	H��2ӡ������fp��ٰ1�/���|���]�����&��3?z����3�9{C���R}�?zZ���i�G*�&����L�1���Ϣ2����.`�՟R�_Gsv~�}�(	ν�,掿�э��2-,�ΠH`�iF��Q�VP��T9ZG�4X�!x� f�?� ~���M��
���ڨ�ƿ�8��ss�A�����<֯� ���f3�.�\o�B 4�����?H�t}%;Fڎ0���8�����1 �`����߉|���A�\��<��,F\���r`Cj��K���Z)v;�����Nz=B��;�����*�|�%蹬ia�f���$
] g୙�Lm��-�(�@��`��	���K7#���
�g1��$i����Wȇ���Ѡ�f搂lo�)�V]��O��f�v�R��<P�C�Q�'<oS{(p�̈́�G�R4L#�<puIH��Ju���;��h�6�E`r3���9�h���傘�4D��.��Tn	4Z���Ԙp��$�T+��E t� b�n�D $�}��h\�H l��-aAlb���9
�~/�	E
k�|�A�^C�i)� ���_?}�����3��,$b~���q�c�����i�w?j�:|�GJ�Ȋ����F��L��SX%(R[x3�|�]N�e��=�4����:��	��\�ϝ�~�5�X3��ĸD�v�1��ۦ{(�	j������R���,���s�M�B���u�;��[��4��dV"Zh63��w���a�ϙ��
7֤� \6|�|��:�d �%��נ�}��e��t�i)`M�9�tbb�,�f[X��"QW
MG�E<������7�e�aҞE����(Z�<F�=��2���T@��̴༙�Q;���t�q��;0�o1G°�8ݣm`%˘1H9`�@��C��ǖ'\bLOR` '�`\D�BIF/�|�ā��NL�ۉBڦ�\��.�N�>�;�cm͑���)Ĵ.�4��Q"�C5��Z��O��4��D��,J���D|s�Q��H�xЦ{��4����E��	��12ftD�Nl:��o��L���W�+�8iS�9�Y"/QC��Ю����ٜ������+Z����m�/i�c�zP��8#�s�0z�,�i�0�գI����I�Ƨg�����Z�^���,�"Q�$t*߯-� ��9į���E��ҹ��ݖu��(�T�ͿG�8���;�ڗ�����d�c��;�Vw�(Hs�%qk\,-��#�52���&R6bP}�����>NXȦ��lD64p�  /1J�gΦL˩}�9U43��&{&��	�A�Mp���1�H"�P&0�;�v��!�d�J@zt*�b��ѷ���9���M�3��/6�WR���S>�S�u�z�4 E��A�WcP��Ĝ;��H���l;/�c�A��-�M���D]Y ����pz(�N�F���Ζ���9���Ki'��A�����a����I�%�N`̦=¤�.P����[B�m;H	�G�DM�	8�sI?'�V��舯��8\��U�eb|zY��Ե)9�[��,]A��
�.��e�| ����l�tƭ�0�0Z�A]���mD�[�'�%�<khx��t��8	�+�ksV���W�T�1P�EP�K���#W�#z#Gk�X�ZB>�����H�/mC7; ��bmk�(lND����b�D�#Q�;��A �*����Cӕt�:G�B��~|e7Q@'�B1W�|�	���݌&	�U�*�(��/���ٌj31�2�2]�Y�힔[ǂ��%&Tڪ�^M}��gM��٦x�)-'k�����y�A�mqΖ�J3�h��
1�r�8���I��3p�2+�F���T�viڠDhT���DX�� J����z8�Y4HM��㱲�s�=g���Y�R��}ߢv�ykrr�������T=��L� H�����m�ZX����5.�K�h�|��壎��A;g4|����д�ܚ�y�\�'���i��w ^��z�v* D���R:��aη4튐7�lO�4m�\�h�4��uV��i�#[{�ˎئ����i͑E`̖vp�.�ɾd��Ѡ�G+�P*nw�m�Mi��F.q�(Vz�WZ0���-��pʺ0�~�5��E6kbA(Mc/X@�&�{b�O�=M�lj���,�U�,�5�ml��q�V
�1�d���\�]m�c\B�����s��j�E�o�0tà+�CpH��)�T��ԤI�R�  �3}pncN�����1�1�Tg"Yj�PfՕm�`nJi�D�9Vve�A�;��ԩ�?���������燿��oz�\U�����C���SK:��_Ҵ��d>6�����Z���X�f�ޟ�3�O�ީ�����������|+Pr��E^~k-�&g�����+7�e�"����C��`Vo"N���{�G���ML��ָ��"KM��%��֊A��AO�u� �|�,mXn���f.f09V���h�Tʰl��Rl1��ڬ���-��Bڋ��2�R���J��v��,���t�1�&G|��$���VAʎ����\�����<k���*u���v��K0�eҷ����kF��]C�ϟ��h�����Y:1�B����Ri7�&�X��U�DUw���y�\^v�e'���Xa�iDr|H�Q'��ulh%�@(�����9U@t�8 ��]0gD���\.ӂ����СC;�y�G�y�����I�m#�!��Ly�u��4<��z����	�ʗv����
�5<y��+V��ٸ��2�J��fS峵t"�fr0�hn-�zZ��]�e)6[ A�En�h�4]Nc���9����2{*�L�J+�V�AQ*�Q�����2L-�BΊO'�w�9m؋�%Q��5\���Y
Pv��Fh+�1�|^'Q.���i0d��T2ca������Ү�.k�6�?�G��Xƿj'�yS���<���Kog����u#�50ո���g�������رI�hB�y��]_kUa)�.�Ll�7��uo��.h6���E��'�S�P��A�/�M@��鎘�S����rƎ����@��&B9��?tV$��믿��fV�X,��FCTg�j�>{�l�~���;�|�7~�7�A����Fୟ��P����8�m�
�^�u�ӵ�&���\V���X'F�e�@M\j���LiM��l	B��Ĭ3�*-�!0�zZ G���Z�ǚ:�bu\5�3ha�����-q�/0�J��:�A):vA����\;�>w��|��� F�f'�	xR@�ӶD��fi��*m�� Jl)¾p�}k��Qd�^��/Ӳ�� 2/�n{�~8��h�*E��!�F=�Flz���4�
3��u�v�̕�tA�����c�Y�C �"<��:�`W����`����yW����O���)F
�ǎ�v�`Ֆ��!̘�-��&�_)��2��H(ѵ^� �F}��a�ƍضm+��>�%�����p��1�9w^(���b*�,{������&e��8�\��(?��O����o�{n�z��G��e^R�3�1�	=��u���D��344$ ݈hTG��	R�RD}Y����LۮX����5.�0�
�J+��rR�����6�I��	kC��g�#�����h��3�X�,��q+g�|�̦�Iu9Y�[��;��hQS���I��X�Li�2c��,�Ŝ �b0�&��G)�98k5���(���D���TM��5c&���)���5�r�n#�3)�T�*�:�D���ij�B1UF��	ag�bG
 �l���lگ03Hmb4�f�ք�c�v��i-��t�0�]}���@Oc�j_D@�hS�*U���g�ϰ�}X����� ��>#��֢~��J2��j+��j��G��i�Xr�����~��x����_����F�ݍ]Z���c�#}Μ�(�J�M��tM�R��5����ڏ?�� 8���������6�n3�x�e�����N`�2�������g�aѾdW|�����ӧOo��|�R��C�r��AQG��[���*5`��P����-k�N������Ӿ��5MM��!�
�ĭq)�κCvd���b	%[���I��4i�Xq���#Ԁ�Lv�U,��������� +D����+mÓ���Y�7�z�!��>f ���ؤ;�#se�+�N�w��f<���
 ��kz+�&<��B�!/}��{����vlI�BT�et���8M5\G�Q+��W��\�xJ�Ԣ���2��u9]�ȝH��LP(��m�X���/*.-��R@A�EX��x#��K%G)��Qh�9�����Ah��*	fQ�=����'b���a޺�&~?
��-T�.M��V��X��T�km6;�KE��~4;Mj�X4c��O�Y�tmjF�#X��15�˓
=<� %���	Qߕ�S@8��.���fh?7;5 P`sl�
�%�܏/v��L�]�@��������7�R�S?lw������]�#�i�V��7��/��^�v�����2*�m�ǿ��_�׿���t?��gP���9�C�f:�O9�@E�-�x�L2f�%���������_�_���a�
�(�ُ����=]�r�7��k��l���=,S���|��{����sk`۶m{hc���-k\o޶�|83`���K�!�9�� �:I�/�r�������n;�j�B�Aj�q�{Y�v�ZwI���j��f]x���/�}G�gdďxԍ���K�7��bN��Q����0�)��AԱ麕C�?wk~ƪ�h�%I��}��5d�3��d'�`���&�Mu�N_œ��P�9"NZ�J���K�2��,l��Ku���EE�m��؜��
J�&�ޟ64:�+E���zJ4��d�PG�0!�.悐����u�Q��6"Bkf�z� X �L��O�����$�1�;B��v��#�oE�E��� lԑ���P)%h<K�hv�*:t��h;���i��V`�8?i+j���Ǻ}�	�;��hh�n��ˬ$P8;9����R�_�(ӵ�5���:Tπ��,�ϰ�bx�j��f����2S�\�3~���,�1�F�L�,V_&�U񾋞�Ҡ�L���^1�4��1�p�{q}�J�3_�:�����e�>bj�l�,�O}���ƿ�׿���S��"�j� C���l�H���k�DjS�n���޿�7�
��ڃ��������y��T�1�c��uL��}����5�V����i(M{s{���ӯ�Җ����D��A�i�).�F�/nEj�Xrwd�O����������+�\/b��饉o�1v@`�gc[��y���Iά���,�ۖ::����j�g9Q�䊛^b�
�ujx��عc�'.f�OC�T���9���,{"��
�������|#<�1�=�d,YE����aB�쓮5{bc�3@ͬ��6��]A�����*u���&<7v�)Q�=0l�_@�Z���a�c� ;o�ۯ��b��gq��ۘ��}�K_E���*��<���ҏ���s��y8��#(����X�	��Î�F���O����[�a��;�����wA^�ӧq�G?F�F�a4i�39,Mك[vb��G�k����a��98^��ށ���蟙�mg%#ú_������i�Ҩ������:�N���s��\��T�'p�/OAڅ`!�����e���s���� i�Y�cG������6�9]���ǲ9��ӌ�w�ʇ�!	Rݷ<�8�X�x��ܯw�}��_�e<H �s��%�}rzG����<fh1P*U0�߇u�G�{�.�U��<EG�䓏�ьq��,N���<rb�v���=�S�+H�$�,�4ڴOS���dA�@�NǸb#swd�j9�����B��y�(�
IXu8M�r��#[�0�iZE䩗G�\V�7䣕�>ϵ�n%�1N��u����'4�ri�P�xQ/֥k�%K;�_/��J��A��Jut�^�<��[�{�?�&2�h�Y��f_�V�h�n	�N*�Y�
u�M��u#�������8zV�a��[00�5�	���[x�I9�ԑ�胷i�h��.M!n5pf�w��i`��ȩ������u�7�ZX��wx;���w����ع[o��! X�	�a��;v�����asz/�`�u�-�X6���``d��V�UG��8*}U��=��a��K�mD��~_���M������q��9�Zl�%i�-�Ў9A�"g)��I�2�A�P�h�	҈n�x�����J��I2�$�CϚ���a ڴ-[��_�
�{�NY���Ë���g�y���&.M��	Ŭ��ƍ���#���f���C��-�~�SE�ò��NRث��Wܠb@H2i�VB�ȇ�8G��b��Ap�+��� �:ȴe[-�"����  y55��1d���텶���8��qJc�K���:UhЋm��D��[t�~i/�,5�'�\t9���'�����Z�lQ����5�_ž�{���'9�g��[�~iƙ�7)�b�^e���fn�
G�y��©��,���x�)*�"֭� e����ޏ��B��o��wފx����p�^���1j�{`MxQ؄ń�t���l�{ѤER���c��_ �}DU�3� "��{H�����~�G��=[7"��>:��!j�' .��I��C����&�t#u����۠�>l��^�O��X8q����{�����TwmCi�(���}3�y~��Ә<~~�����i. ��u�h~B�Cu�vl�m/��F}�μ�ֹjq �nu`[��o�R2��&ٷ?]�^1�F�
��<G V��ᡇ�SO=!
3��i�}��g���8n�N�/�HB�����\���,�=���:��<�����~����Գ~�'w1g����x1��o���6�	+ݜ�����[��~��|rw=�XH}�`y�������ک�|�R�
D�cѹ�/��^ui�����21�Z���h
ik���o���aЊ��ն��"�y�%��4�nX7��K��ݷ���CG�㍷�՞I���ݛ]��Z߻	�HESĹ�v�da��I�~�L��B��Z��0u$��19�;�ߏ/%���ı��P�̠�F)�c��<��zK=��0�y�z׽��Dc3b^uhX �4N׬M�c`�n��Ѓ�D+����N��F�����D��TO��8(��/ �~�0J{v�41��%WMF����Q��}+��¦Z����64�[>�0���� ��P=ƶ#�����l�b�<L ��i�0z������n�Eڱ:yI�F�����T��
#�Dͺ�o�nVg�r����R��sM8�GSCl\��{�qE	#S�/�������̹1jW��-�����`�r(�<�[-��Z��il۶�O�����*
��`$�9Ntd��l(�|��`�Q�XIr%�H�gsj�nVq�q���؋q�ǦSBG�눉D��C���Z�:_�|PX�0���j���6�yT��J�\��K���5NI��~-�Q��ע���6)'��,{떍غiP~���R���\�Tq�0@(.��r���]Wyd�2��Ku�9@Y�9*Wi��E`�����d���~�߽ع8{}� ��<Ͼ��׆a��nqGh1�y�-�&���-�+�XkϡMߋ�܆m_�2]���7_����X�S����0����{�ƆM�Tq��e�v?7Z��#��q>�X�C�O
Et@1,�D7���9�wT������*P"@:1��w�af��������P�h}�T�:Fx��_���z��kڗ��8�Pd��������������η�r�T6skr-Ձ�!�e!*^Y��GCZ�h���z"�d��|��l݄}���Wl8?6���Y=~���.kw�p�
���Z�-3��㹋c�xiB��t�Y����lD �^�_In���~~�c��	l0�.K�{��?I�0M��~�q	�>A�A��'I�(�JPɬy��A���bM��.��H5�D#�1ߍkx�U���*��FQ�!�.�Mg�Dj@H��4������T�������������M2�TQ5�4F]3�e@���Y��oF$����FU�?/]����L��K0�S� -1z�Nl� �r��~�΅��;x��[(}������î2M��0��3-�~p��h@;{�X�n}���-��_��CG��-@��V�`�ԇ��38��������}`��_J�3?�kr�(k_�/��U��u��  �ϵ�䖵p�M_'�Gqf���anb�sah�u�q����W^C�8K��[��|���� j�O`s_�ީ%����*�>ظ�0��G�E��oUG��ּ�`cm�����+1ج�RM������n{��r�$ �U�2�CCè�j[�w��LL�ȢS�a�*�)Ȣ�(.5�X�a��Kz�Jh��r�(Q��Sn)QDo��,Q�qs�v�b�޺���W�����j}��u�W�]%q�A8n�瑔�ߙN���-l�zS��S)t��Sqt�.[}^�\���fv��a��ľ&�<B+W�A��R�����L�q:��f��y���iG\Ι���P�7E/�pS��(h!�;�݂�Գ���u�w���d VFa�t�	�tu��47T�x�D��L�a+-sh"���TTJ(ܺ��U`�V�pN��*A��r�vm�_�E4��|�s?��~;.����ݷ��ؓ4���B�:>�������ˣ�q�ã�p+G)`�=������I�O�Ʊ��>���ß�<�z���#ʵ:���j��[� �#��0%�@���CY��QIT2�G;Ql�����K�Wh�C�6��6
x�;}�0��6ѳ@�%@�/�g�Aؙz�bZ���c~��C��<�����_ϡ0�@ډ5�T�6ܼHiso���+	)�FMC��/�m�헱�S�+8{�<Μ9O�nS���� 8��9���`p&@��Q�4$�lY�f[�me>��є���<�[�b��$��`�-Bu���ʃiXz�B�4H�z�T�ۋ3V�8��A {�tͬK�H���� �iG���V��;q�I,�]��(%ؗc�b�I'S��[�7x�<��|*N�]��,x����,��*b0M�����2���	��8��ѣ�R*!�iB�����P.ѡ	5 ���(Xe��1�	�pNG�'e�L̠���*���~�v�V)�b�.K�dT���ڈq��T�;���_�må7��k�ӸΠ��$�sǝ��
q��	,l����`�Jd᥋cH^�):��k���}C`zh�z�i8+V����~N�ņ�!<}���������G�RSZ��(±�ꥧ�i@�`p� e��+��B	e�H"xQ��P�~���D�Lן�����۸�.��WFe�:N��LŘ�G���:��3���|�5$��,�8�ν������w�ҋi^'q�:�,��n���+݁�M�J� �%��%pEߓ��º�0����qz7Z����`����̵��&�EWq����H�߰��.B���Z		T3��J�a2��N����O�\�h4�-0c�i҅��F��~����qk���R�|���!�Q;0�<�A�u��+�*�Kc˗�N�J^G^�3ӓ�D`As�&�F���s����R^.���L6��?z�D�<:���NB��8��sH�f}�@��E�[��������~��#��JRV��?!����kS���W%	V���5�hq9���	�-��g�_����<=�5Z�`�3wa�W��u7�z��0�M;nÖm;q�ݗ���;Q��P�Ǳ�^��i3P��'Q��#"�3q�(aaZ��K�g��m��?~��0ڭXw��7`����U-l��_6n���/�c���$O���t}�oF�0J<6ACr�G�v�ʏ}��[P?sq_  �N{�Zto�BZ(�dәC؜C)�`��V�1���)Tno������� ���	`���k/��! �}��B�WD#L���(�� �O_���
�;�*eT���b�8���Nh��X�j���'r���z��邓T���9��dV�f �f`͚,�$�%�V8Ҝ�ΓX���D�i��rMhk6�W�\A�$����ɟ���I�8�� �:[C��b-1i~T�b-�t�0��A���[�֭�����R�-��o�e3�j� 5 .k���]�P�z����Drw=$���W*	���3QL2�Yj Vy/�J�k|���ɛhe�fIW�z䣉����A�+Xz6�6m�#�ދ�/J�Z+��Ý��R��~�	���da��c'����9nvI,��C�tZ6~ǭT%\/�!��e�6`�6�u$����� �n'�:wo�����3������]��b��A��(�����ڴ�J��6�����1z.e�	�Y�Y�!��؅�Xv/��Q����R%Y�c�;�E� P��P��
�q��V�|W��"�;A�l��c������}3��/y�C�0�+_��o���[���ģ���������}�{��(`3]H�Y����Q�c_��ã����1u��9 ���J���--t���b]���I;��I��c�ʸ*$�<Џ��~4���8M�C����rY��PXNE��P<�,a�s+c��Zs�;�J�c���5[�r�]t����þ�j�l6�ubE�S�y���S�J�Tj[��揥|J��h0�_o��c����Ǜ�x���3477� =���X+W��<����f��X��\�jͲ�����6���S�P�A�u�ԥ�a�	��)2UL�N�V��5�	M�l��z#��G�GQ�Y��TS��X4�-:7O�%��iY��<Yp���L����<�lʊirp�A>����ʱ�<G�����H���6��aS��pnu?2�l)Y�f8�����O�A��;�&e�L��D ��xNN�`+����ob�����afƧ0�"��Kp�m�^A%�/x����'l�`��g�:���fq� Z��gl��i���ǖw���~����4�.��i�/;��j60w�(3�E��:����ՑԚ���� m&��X�8�?�����B�[' PH;�������?���	���Ϝ(���4���L�#
��*�Q�rP�+b��������������c��Ixg'QqS1Y7�D�q���]��OEu/�֢U�D��Y�9�8Z���ӧ�t���;�a��-x��qo-�bq{`�'ױ�Kb�Oe��}�w	���Ry��o�-	:3AK,K5�+������$v���W�g������_��ַ���^�t�g	�m�gU��s꺮=11Q"�V�O�h�X�7#�1g�}��s0���rEv��]Q�p���m�.��DG�$�5�S��9S J�i���#K��D�c��$����YSjw83��6��^ g˄����z�� Y����,�\�1NV��`d�q�|�#͎��$M�}ff����jѤ��*1��M��jOk�����̓�"u�?Xb����=wNRJq[ԙ�Hes�T����Hq3�'(�*�%��<v!M��U��a�VM��C;�|�kb:�;G��Ա����L<��#���G��J�!��cr��;�	9(4�HN�D��B�Zgj����B��[r�%'D��1u�mQE6!$/���UJL���9��Q�^�+�i�u���P�;�Vˊ�J��1&�=������D��d�t��p�Tę�b��]CQr��Eˉ��h3�G�*����"�N�Z���}{w��;����h�/G3EL���pr?/һ��CY����$�6�Z���j�<��0�X�npJW�J�R+L~��_��_��}���]�Rq	t���m��l�����S����C��.:d�@�c̥Y�>�$�}�&O�?�5q7�x��( d��v,&�Ԥ[t��-Щ�X��]�#�Q��Wur��t���݋�Ӆ쮁��b_�6��J����j5Z����s�=�#G!	:4hD��۶y3~�����L%G��;���~W̩<���G����)�R�Feb2_d@�*ϝ*��^���]A��?E����&�X�bz��]�Z�M�0wq}�*����4U]6o�1	G��;��ZBs�+Q��^?5K@B��沔&wWL��/kbB���2�@�EϥA@�!��<X|���X�i�=E��'Q��T��3�f��$��^C?mw��&��#�k��tG/�O�)XE�gX?2�Z}�xt�,~*>�r�i[��e��E�EU+��^r��;F�tӹ�~�J�Şj�Q&T6����O����	���x�����;S������ѓx��Q	�������s���c+%��is�~�e6n��Gq�ܘ�?��˄�<f��m�+PX�|�⣂(�������W���u�����7�x��s��=����7Ýt_��yW��}�$ȁ��ѧFu������rwݤ7���N����K�+���rYɚ׮����.��
Nh!�'
��h�QJ��V��
ؖ�������`�h�a-N���8�����(����'B+Gatwluƙ�9�w�(�TE3A">��0tb�me�|�q��Ħ��}���J�JÙ|�����^l@�����MJ L�v�,k=�^Cr���r������\CH\�0�b�K��$n*T<1�b��9�Rn4|�.�nѱi�cGdj��o�W'a��N�� is&�����Ӊ�	����(J�lu�#l������Y���x��A$}!&��ђ�����JT�j����i�8����!եT��C}�2l�a��:O@�i6j�����1�n��&Ό)��:��r¼��q�����=�߾�s`�D��;�FB���/���-Y<xn��153/TI�N����ϚS��Q�����������{�-�o��[|�?���%I|/���t!��+,��͎�+c��3�/��PX[G?���u|||�������ɓ�����G��[k��b������]�GX>�8���A,{,��P��h9A��)V�� �:H�3��hԮ"����������-�ϱ�48�|�f�������l�C��cL��Z|j�T�D�ؿO��$��8Y:����Ջ�^�1u[j������zG��q��:�����8x��i�w�����7?k]�84��e��t�R+�Ä���L��1H�1����)D�Z���y
�ii�\�8����	�>���
N�V@�ӂ]tqN�zz _ҼC��b�|� K �V#ǉL�����X~E���L�x�]Y(g����}Q��mdNGά��(�%��}r�����3X�6Wa����M��`���v$��&�RA���r����v�<��k2ѬYT�=��B���H�*��+R9p���x��l��eЪǸ�U�-��T�9P;��^|�}�������^�S��;S��_������K/���w0?3+�F~P�R��o�=wߋ'�|wܾCH���X�������y},aP`� �Zj��L�F�~����*V�|���nk4w��;��;p�����ǇL�X�yr�;�BA3�%��?�,�7)���]F�������Z�o�`��M������?��?�J��]'��۱�P�D�鉊�r��,�9E%��L��Bi讵��d\k��uS�t_�V(��cː�f&[�,�+`-z5rem`�a�l�~k����ϑ�
Ӑp��<GK;�[:�������"�"?&��hՕ8T[��@g��h�,��[\Z]�ק_�]_�w,�o�q��8�ҽ�^����/v�e����������N\ ���+����,[�����/�_����c���ϳh��u���!��Zʮ�pW�v3�8�Q��]�*K!�dZh�	��.�����]���~����o���.�u�~�:u'���y\�~=v�؉�[��Ttո�����}mG�g�E��Ńh�Ѓ�=���q�q��7���9s#�����X����� Z�{�j����OE��	u��:�L��?�rO.?IX�QQ��͔
�z�2�dA��n%���M�+A�&�t9�c{�˲�Ltˊ��_No��=�}����<L��G��*�@�
`�@�&ˇ���ۣ�P2%gD0�l��y���D�	^�ND�3-��.�Z��'%r�CM8�g���n�ي��K/c�Z~����g�~�����߇{8�9K��h9u_��i�^����p����ζ�i�i'��/�,�V��X�H.7Drw���}_�}�*���
z��>L�FQ�Z�c�i��q�6�|Rk�.�P&tY�!G�-��/Fo�p�e�����\�bjy�'/�����o����j�Դ�RɶN�L��.�O*@L��Dio�� ?��~P�x�Z��^�����\
���0J���#=nF0�L�D*Ƣ	wlO�Y6J���_|�.]��z�=��o�$�0���q��d i�跙�?}ϼ�^x�U�>yJ����Ծ���#բM-�/ve�D.��X�A���$��A@��C>�^oV�z�Nԟ�(8�2��j0M *�1���[�&�,3 �8�4���7O���j~�y�J�޵^e�)
B?�`rr�������N(�BsLF�g�z6z�L6pV>s&@d�n0=�A�5��˪*�Y��O4p�cs�2��-a*C����*D"  VIDAT�K/�^^��l��9��y8|w�u'v��&f���!�?d��z$`�̙38t��;rG	�����
E��"�N$`�S$bݾ|�T^��+N��*��'/9��Xv�V;�j�XM½(�DL� ��Rē�BW�]��J���lt���)<'���5ȋ3~!�Gdu��St��GL������e��;�s�-�OU�Y]��r��Z2Ѽv���,�Q�=ە%ѯN�rY�"�`�7*jY־�gʩ�,H��SK�Uwc���&�xE����������P�T�m͚Y1'$��qƀ��L���-T�.�}�ޔ`�T�`�8h�̀�U�����5(9������'q۳$u�A�)�V>bn5���P&P`k�׵�=��k--�4U���`(M\�Dd@��qV��\#��x�]�D�Wj�=`ē s1A&��h<����K-����62`]E1��h�f���8�3�~���+��?c����T%�OM�l��MBeD�P2�D�K%wl�>t��ri";�o�;&fk8~��c���+��r��|�Ǵ0L�}O�9��#��P�Yè�q��b�믰��ĭA�A�u�T�Sۢ�J-mN�D�i7���i���"`�K3�6���E�Q��r��R�N�G˲����z���^��	p9Ha�V�e
�e�IYx�WI�=���Q	șE^��yy1x�6�J3Yڄn) ){q��<��ͩ�U6�ս���y��JeBe����f����Ux�����za��/�&����Ğ�@yK�PB�U��p��_̢	Ӻش +���g��a@��P'���x��n�I[��o�nj|�W��.���DsY����� �vx	j�ё�1�|���C�}:�oG�:��Kd`2��k)��aC�$$��u�B9Q�Z6�J��qw7�si �4S!�≶/^V�$Ѿl��fF3^Q�y2a~;ڍ�d왣L�k]��3�*���a�Y[��'!'�z5dx��㜙Lh��,�QN�����Wwk�oY��a�e^��R���):���wa�Kj����ⱓ3}p_s%B5��n���ʘ�
}�Z2QG�^�:�ۙh�|��&o����g����6�r�o$��I�D��-�" �;rMN�ŋ.���<};�%g�%�OCrw��y3�'��`.�)�Ki�W	;q�vt���X�Zily��)��$�Sj�]�2��]���F+���}�L�*�N����N����i�/%C��B'8��ݼJ�|�!�
�t7��	�V�tW���ƫ�T���h�8�j�_�>X���Ƽ��*�g8N����<Yd��k��<��#6#0�%�m��������\\�x�����
���˼���\D +d���Ǩ�����.W�l�����L�w� ]���ofT�����%%�K�����w��P#�(�X�F26�*��g�(sj.kPrwd�W~e��_J_���i�
*��-�ݺ�&9~�>Z��}Q*�Br��uFBUA���:~ڻ|����};��8��J�cG����RLؗ��?���u��%�K���=����U`r��L�e�,�+U�`���nux���g�yu��8�[|0�l+�0^`�J��M�5�oK掴�r��l�}l��N�#�|4I9�cp�Y떙�Ds�˥ .�>�Z�����T�"ʥ>)�h��pz�T9&���� ʰ��*��nE�O���6�bQG6�]��F+��i��u���s�q�\�Hu^\�iw��\r������(�4��d�ß9��ą ����J�>"0&5�@�l$d��7v(3���4y%�v����GFز$���k�S,s2�������?K�o�d�\W���Iήb,�:I(���h�"��+y�J��@��m��%/�ru�Z����RG���*7����&�jz��U�\��:�Ǌ�6�ht?�^R;�Rc��`Ρ�y�CCO�#�Z�W���XYrY[���5.'�́�N���h�Dcž%�sGB%Nf��z�HȂ�(h�s��]�ϱ�&a W�P]����|�,�ݕن#�b�������lÿ!��?��۞�V|e�5-'ֲ��r�e���H�K8@�A��J^�P��"���ȸ#>��Zh�Lf��ʯ��v�R�Ғ}�,�����d�q�Z�T���v���4��X)�6�M�A������K�R�/��fy����^e�R�0J9��J9#51f�%�1_�m�����Gq��wbn�)�P�����r�B��s�<�P�$������t��TI�Ch���cs�A�ϣ�~W\C[�"��Һ�=@.�\����ha���ӡ���K����-�]�틶[��i_/VSW/+ΕBKC���pۆ\;[?6��O*�����صs+��%�s��TΜ���U+gP��S�ĭq�A����GN:�8�ɏ5Ga�E`�$�M\v��������<��əH`�T�⩧����M��.8dt��Z������L-�	��u���x�O��	�lY��e��觶-�v�Ӿy^��cr��j�I}I?ǫýNwzU�-O~6G���E��u}P�\������[{�5�Jj�+��ڙs��>^�:��R�n�W�Q,�T|X9��\�F%qk\�v\�PRL��X�O�\�S,K�rV~(j@ԃ�	�_A��:L1�Qd1M�V[�^�V��Fq'��+kMt(��Qv�Djq����s�ހ�}��^2���1�H�5�*�eR�|�v�w����y��J^ѫoGJD�%��9��C���N�P̯JϦ��)Ό�b���+�D�'�?K$�6�2������R��I(c	SEq����_�k�֨� n��ǎ;��
:͖T)Ta� Ǖq�̈́L�!�(2
/�pp���f����e<H�:��>x�M�xߴH���� �i��w=�rO�qdŁ�#$I[�������+�S�Sr9M���+.К�y�z� �����%vRߌD;�
!��y߭��/�3&._���s���_6��������d:#��2��#��Z�o���D"����ʁ��|j���5.�⍜�
*��0B�\�4S�V}}}�*';XYj���#R#�*���W�6�˖�M,�?�%�I�],��\�c��//�r%�"4�p��R�.�Of�Ɍ8�7���xr���f~[N�5扙��
��T*� nJ�ָD�ی�x��7����ʎͪ��\r�%��)����t�A�ө#�5'9�[�R���>��j�<�Q����Bs�Pa%�%�\r�e�	/�ٟ����F.kNr��ejjj�ԩ�o������^q(��>�qtq��aj[;M9+I2����Ye'V7�����߹�崒f�1i[�j�'[��̹���V����u��d���R�Υ:�p�Dvj���$s��;G���}8�H��cx;_z}ni#K݌���n�P۩6���o�n�^z��n_�>���^��,!�����=Y�6ǒ6���W:�J翼�ׇUu�k�_��K��A��<�=/�,���~�g��?�T����:�������|H�O�*U��U&
]�|�>�,�d�����nCf�YZ���r2�x<2�9ƌMV���c��L��}.qs��K'w�Dꤰ[~��^*�O�Wq�6��-9�^}��>�6��='�jՂ 8933s��9�A��T�������h���߹�K.���W �4���>~���g��1�R��$q��� �gr�%�\r���,��x��ٹ� .�\r�%�\r�e5J�r�%�\r�%�\V�� .�\r�%�\r�eJ�r�%�\r�%�\V�� .�\r�%�\r�eJ�r�%�\r�%�\V�� .�\r�%�\r�eJ�r�%�\r�%�\V�� .�\r�%�\r�eJ�r�%�\r�%�\V�����j-�rW    IEND�B`�PK 
     ��/Z.��\n) n)                  cirkitFile.jsonPK 
     ��/Z                        �) jsons/PK 
     ��/ZA���/  �/               �) jsons/user_defined.jsonPK 
     ��/Z                        �Y images/PK 
     ��/Z�ȅNܶ ܶ /             Z images/d20a931f-9d34-4029-b213-4c0e689ce6a6.pngPK 
     ��/Zy����� �� /             4 images/cd711d72-4439-4fb4-bf4b-39cbaf4dbd75.pngPK 
     ��/Z	��} } /             � images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     ��/Zd��   �   /             v-	 images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     ��/Z#���5 �5 /             NN	 images/4ae07c11-480c-44ae-b2c6-f8186e930d96.pngPK 
     ��/Z��5�) ) /             |� images/fbc1041b-f35a-4c82-8c92-5608856c8a22.pngPK 
     ��/Z��d[�  [�  /             � images/42ade947-84bd-4266-8f8d-47ba602ec33e.pngPK 
     ��/Z�I��5.  5.  /             �K images/ec55ee1b-9bfc-4adc-bb90-2198f3917cd5.pngPK 
     ��/Z�J�?& ?& /             z images/fae5eb44-bbe2-4b21-a13f-fb7a66868d1d.pngPK 
     ��/Zp&ر  �  /             �� images/aaaf988e-4d8d-46a5-ae55-a0506af48a51.pngPK 
     ��/Z��[.�	  �	  /             �� images/e8fbe2d9-26e0-4ccf-9f9e-bb43371c63c2.pngPK 
     ��/Z��`  `  /             �� images/95d79837-2dff-4c75-b12d-e13dc3081ed5.pngPK 
     ��/Z�l: : /             b� images/bce349f0-9fdd-490b-ade4-f6d95f909232.pngPK 
     ��/Zִ$�� � /             �� images/4fd5fc97-bc4f-4740-9bc3-7af0136a9299.pngPK        �   